`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module RetimeWrapper(
  input   clock,
  input   reset,
  input   io_in,
  output  io_out
);
  wire  sr_out;
  wire  sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module SRFF_sp(
  input   clock,
  input   reset,
  input   io_input_set,
  input   io_input_reset,
  input   io_input_asyn_reset,
  output  io_output_data
);
  reg  _T_8;
  reg [31:0] _RAND_0;
  wire  _T_12;
  wire  _T_13;
  wire  _T_14;
  wire  _T_16;
  assign _T_12 = io_input_reset ? 1'h0 : _T_8;
  assign _T_13 = io_input_set ? 1'h1 : _T_12;
  assign _T_14 = io_input_asyn_reset ? 1'h0 : _T_13;
  assign _T_16 = io_input_asyn_reset ? 1'h0 : _T_8;
  assign io_output_data = _T_16;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_8 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_8 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_8 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_8 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_8 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module FF(
  input         clock,
  input         reset,
  input  [31:0] io_input_0_data,
  input  [31:0] io_input_0_init,
  input         io_input_0_reset,
  output [31:0] io_output_data
);
  reg [31:0] ff;
  reg [31:0] _RAND_0;
  wire [31:0] _T_8;
  wire [31:0] _T_9;
  assign _T_8 = io_input_0_reset ? io_input_0_init : io_input_0_data;
  assign _T_9 = io_input_0_reset ? io_input_0_init : ff;
  assign io_output_data = _T_9;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= io_input_0_init;
    end else begin
      if (io_input_0_reset) begin
        ff <= io_input_0_init;
      end else begin
        ff <= io_input_0_data;
      end
    end
  end
endmodule
module Innerpipe(
  input   clock,
  input   reset,
  input   io_input_enable,
  input   io_input_ctr_done,
  input   io_input_rst,
  output  io_output_done,
  output  io_output_ctr_inc
);
  wire  SRFF_sp_clock;
  wire  SRFF_sp_reset;
  wire  SRFF_sp_io_input_set;
  wire  SRFF_sp_io_input_reset;
  wire  SRFF_sp_io_input_asyn_reset;
  wire  SRFF_sp_io_output_data;
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire  _T_19;
  wire  _T_20;
  wire  _T_22;
  wire  _T_24;
  wire  _T_25;
  wire  _T_26;
  wire  _T_28;
  wire  _T_31;
  wire  _T_32;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_39;
  wire [1:0] _T_45;
  wire [1:0] _T_48;
  wire [1:0] _GEN_0;
  wire  _T_50;
  wire  _T_53;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_57;
  wire  _T_58;
  wire  _T_59;
  wire  _T_60;
  wire  _GEN_3;
  wire  _T_76;
  wire  _T_84;
  wire [32:0] _T_92;
  wire [31:0] _T_93;
  wire [31:0] _T_94;
  wire [31:0] _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire [31:0] _GEN_13;
  wire  _GEN_14;
  wire  _GEN_16;
  wire [31:0] _GEN_17;
  wire  _T_97;
  wire  _T_98;
  wire  _GEN_18;
  wire  _GEN_20;
  wire [31:0] _GEN_21;
  SRFF_sp SRFF_sp (
    .clock(SRFF_sp_clock),
    .reset(SRFF_sp_reset),
    .io_input_set(SRFF_sp_io_input_set),
    .io_input_reset(SRFF_sp_io_input_reset),
    .io_input_asyn_reset(SRFF_sp_io_input_asyn_reset),
    .io_output_data(SRFF_sp_io_output_data)
  );
  FF FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_19 = ~ io_input_enable;
  assign _T_20 = _T_19 | io_input_rst;
  assign _T_22 = FF_io_output_data != 32'h3;
  assign _T_24 = FF_io_output_data != 32'h1;
  assign _T_25 = _T_22 & _T_24;
  assign _T_26 = _T_20 | _T_25;
  assign _T_28 = FF_io_output_data != 32'h2;
  assign _T_31 = _T_28 & _T_24;
  assign _T_32 = _T_31 | SRFF_sp_io_output_data;
  assign _T_39 = FF_io_output_data == 32'h1;
  assign _T_45 = io_input_ctr_done ? 2'h3 : 2'h2;
  assign _T_48 = io_input_ctr_done ? 2'h3 : 2'h1;
  assign _GEN_0 = _T_26 ? _T_48 : _T_45;
  assign _T_50 = FF_io_output_data == 32'h2;
  assign _T_53 = _T_28 | SRFF_sp_io_output_data;
  assign _T_58 = _T_57 | io_input_rst;
  assign _T_59 = ~ _T_58;
  assign _T_60 = io_input_enable & _T_59;
  assign _GEN_3 = io_input_ctr_done ? 1'h0 : _T_60;
  assign _T_76 = FF_io_output_data == 32'h3;
  assign _T_84 = FF_io_output_data >= 32'h4;
  assign _T_92 = FF_io_output_data + 32'h1;
  assign _T_93 = _T_92[31:0];
  assign _T_94 = _T_84 ? 32'h2 : _T_93;
  assign _GEN_9 = _T_76 ? 32'h2 : _T_94;
  assign _GEN_10 = _T_50 ? _GEN_3 : 1'h0;
  assign _GEN_11 = _T_50 ? io_input_ctr_done : 1'h0;
  assign _GEN_13 = _T_50 ? {{30'd0}, _T_45} : _GEN_9;
  assign _GEN_14 = _T_39 ? 1'h0 : _GEN_11;
  assign _GEN_16 = _T_39 ? 1'h0 : _GEN_10;
  assign _GEN_17 = _T_39 ? {{30'd0}, _GEN_0} : _GEN_13;
  assign _T_97 = _T_50 & io_input_ctr_done;
  assign _T_98 = io_input_ctr_done | _T_97;
  assign _GEN_18 = io_input_enable ? _GEN_14 : _T_98;
  assign _GEN_20 = io_input_enable ? _GEN_16 : 1'h0;
  assign _GEN_21 = io_input_enable ? _GEN_17 : 32'h2;
  assign io_output_done = _GEN_18;
  assign io_output_ctr_inc = _GEN_20;
  assign SRFF_sp_io_input_set = io_input_rst;
  assign SRFF_sp_io_input_reset = io_input_enable;
  assign SRFF_sp_io_input_asyn_reset = io_input_enable;
  assign SRFF_sp_clock = clock;
  assign SRFF_sp_reset = reset;
  assign FF_io_input_0_data = _GEN_21;
  assign FF_io_input_0_init = 32'h2;
  assign FF_io_input_0_reset = 1'h0;
  assign FF_clock = clock;
  assign FF_reset = reset;
  assign RetimeWrapper_io_in = _T_32;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign RetimeWrapper_1_io_in = _T_53;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_57 = RetimeWrapper_1_io_out;
endmodule
module SingleCounter(
  input   clock,
  input   reset,
  input   io_input_reset,
  output  io_output_done
);
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire [31:0] _T_20;
  wire [32:0] _T_22;
  wire [31:0] _T_23;
  wire [31:0] _T_24;
  wire  _T_28;
  wire [31:0] _T_39;
  wire [31:0] _T_42;
  wire [31:0] _T_43;
  wire [31:0] _T_44;
  FF FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  assign _T_20 = $signed(FF_io_output_data);
  assign _T_22 = $signed(_T_20) + $signed(32'sh1);
  assign _T_23 = _T_22[31:0];
  assign _T_24 = $signed(_T_23);
  assign _T_28 = $signed(_T_24) >= $signed(32'sh6);
  assign _T_39 = $unsigned(_T_20);
  assign _T_42 = $unsigned(_T_24);
  assign _T_43 = _T_28 ? _T_39 : _T_42;
  assign _T_44 = io_input_reset ? 32'h0 : _T_43;
  assign io_output_done = _T_28;
  assign FF_io_input_0_data = _T_44;
  assign FF_io_input_0_init = 32'h0;
  assign FF_io_input_0_reset = io_input_reset;
  assign FF_clock = clock;
  assign FF_reset = reset;
endmodule
module AccelTop(
  input         clock,
  input         reset,
  input         io_enable,
  output        io_done,
  input  [63:0] io_argIns_0,
  input  [63:0] io_argIns_1,
  output        io_argOuts_0_valid,
  output [63:0] io_argOuts_0_bits
);
  wire [63:0] x332_data_options_0;
  wire  x332_en_options_0;
  wire  RootController_done;
  wire  RootController_en;
  wire  RootController_resetter;
  wire  RootController_datapath_en;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  retime_released;
  wire [31:0] x333_number;
  wire [31:0] x334_number;
  wire [31:0] x335_number;
  wire  RootController_sm_clock;
  wire  RootController_sm_reset;
  wire  RootController_sm_io_input_enable;
  wire  RootController_sm_io_input_ctr_done;
  wire  RootController_sm_io_input_rst;
  wire  RootController_sm_io_output_done;
  wire  RootController_sm_io_output_ctr_inc;
  wire  _T_477;
  wire  _T_479;
  wire  _T_480;
  reg  _T_483;
  reg [31:0] _RAND_0;
  wire  _T_489;
  wire  _T_491;
  wire  _T_492;
  wire  _T_495;
  reg  _T_498;
  reg [31:0] _RAND_1;
  wire  _T_504;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_508;
  wire  _T_510;
  wire  _T_514;
  wire  _T_515;
  wire  RetimeWrapper_2_clock;
  wire  RetimeWrapper_2_reset;
  wire  RetimeWrapper_2_io_in;
  wire  RetimeWrapper_2_io_out;
  wire  _T_520;
  wire  retime_counter_clock;
  wire  retime_counter_reset;
  wire  retime_counter_io_input_reset;
  wire  retime_counter_io_output_done;
  wire  RetimeWrapper_3_clock;
  wire  RetimeWrapper_3_reset;
  wire  RetimeWrapper_3_io_in;
  wire  RetimeWrapper_3_io_out;
  wire  _T_529;
  wire [32:0] _T_532_number;
  wire [32:0] _T_534_number;
  wire [32:0] _T_536_number;
  wire [32:0] _T_544;
  wire  _T_547;
  wire [32:0] _T_549;
  wire [32:0] _T_557;
  wire  _T_560;
  wire [32:0] _T_562;
  wire [33:0] _T_563;
  wire [32:0] _T_564;
  wire [31:0] _T_566_number;
  wire [31:0] _T_580;
  wire [31:0] _T_584;
  wire  _T_585;
  wire [31:0] _T_589;
  wire [63:0] _T_590;
  wire  done_latch_clock;
  wire  done_latch_reset;
  wire  done_latch_io_input_set;
  wire  done_latch_io_input_reset;
  wire  done_latch_io_input_asyn_reset;
  wire  done_latch_io_output_data;
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  Innerpipe RootController_sm (
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_input_enable(RootController_sm_io_input_enable),
    .io_input_ctr_done(RootController_sm_io_input_ctr_done),
    .io_input_rst(RootController_sm_io_input_rst),
    .io_output_done(RootController_sm_io_output_done),
    .io_output_ctr_inc(RootController_sm_io_output_ctr_inc)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 (
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  SingleCounter retime_counter (
    .clock(retime_counter_clock),
    .reset(retime_counter_reset),
    .io_input_reset(retime_counter_io_input_reset),
    .io_output_done(retime_counter_io_output_done)
  );
  RetimeWrapper RetimeWrapper_3 (
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  SRFF_sp done_latch (
    .clock(done_latch_clock),
    .reset(done_latch_reset),
    .io_input_set(done_latch_io_input_set),
    .io_input_reset(done_latch_io_input_reset),
    .io_input_asyn_reset(done_latch_io_input_asyn_reset),
    .io_output_data(done_latch_io_output_data)
  );
  assign _T_477 = RootController_en & retime_released;
  assign _T_479 = retime_released ? RootController_sm_io_output_done : 1'h0;
  assign _T_480 = ~ _T_479;
  assign _T_489 = _T_479 & _T_483;
  assign _T_491 = ~ RootController_done;
  assign _T_492 = RootController_sm_io_output_ctr_inc & _T_491;
  assign _T_495 = ~ RootController_sm_io_output_ctr_inc;
  assign _T_504 = RootController_sm_io_output_ctr_inc & _T_498;
  assign _T_510 = retime_released ? _T_508 : 1'h0;
  assign _T_514 = io_done == 1'h0;
  assign _T_515 = io_enable & _T_514;
  assign _T_547 = x333_number[31];
  assign _T_549 = {_T_547,x333_number};
  assign _T_560 = x334_number[31];
  assign _T_562 = {_T_560,x334_number};
  assign _T_563 = _T_534_number + _T_536_number;
  assign _T_564 = _T_563[32:0];
  assign _T_584 = _T_532_number[31:0];
  assign _T_585 = x335_number[31];
  assign _T_589 = _T_585 ? 32'hffffffff : 32'h0;
  assign _T_590 = {_T_589,x335_number};
  assign io_done = done_latch_io_output_data;
  assign io_argOuts_0_valid = x332_en_options_0;
  assign io_argOuts_0_bits = x332_data_options_0;
  assign x332_data_options_0 = _T_590;
  assign x332_en_options_0 = RootController_datapath_en;
  assign RootController_done = _T_489;
  assign RootController_en = _T_515;
  assign RootController_resetter = _T_520;
  assign RootController_datapath_en = _T_492;
  assign RetimeWrapper_io_in = 1'h0;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign retime_released = _T_529;
  assign x333_number = io_argIns_0[31:0];
  assign x334_number = io_argIns_1[31:0];
  assign x335_number = _T_566_number;
  assign RootController_sm_io_input_enable = _T_477;
  assign RootController_sm_io_input_ctr_done = _T_510;
  assign RootController_sm_io_input_rst = RootController_resetter;
  assign RootController_sm_clock = clock;
  assign RootController_sm_reset = reset;
  assign RetimeWrapper_1_io_in = _T_504;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_508 = RetimeWrapper_1_io_out;
  assign RetimeWrapper_2_io_in = reset;
  assign RetimeWrapper_2_clock = clock;
  assign RetimeWrapper_2_reset = reset;
  assign _T_520 = RetimeWrapper_2_io_out;
  assign retime_counter_io_input_reset = reset;
  assign retime_counter_clock = clock;
  assign retime_counter_reset = reset;
  assign RetimeWrapper_3_io_in = retime_counter_io_output_done;
  assign RetimeWrapper_3_clock = clock;
  assign RetimeWrapper_3_reset = reset;
  assign _T_529 = RetimeWrapper_3_io_out;
  assign _T_532_number = _T_564;
  assign _T_534_number = _T_544;
  assign _T_536_number = _T_557;
  assign _T_544 = _T_549;
  assign _T_557 = _T_562;
  assign _T_566_number = _T_580;
  assign _T_580 = _T_584;
  assign done_latch_io_input_set = RootController_done;
  assign done_latch_io_input_reset = RootController_resetter;
  assign done_latch_io_input_asyn_reset = RootController_resetter;
  assign done_latch_clock = clock;
  assign done_latch_reset = reset;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_483 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_498 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_483 <= 1'h0;
    end else begin
      _T_483 <= _T_480;
    end
    if (reset) begin
      _T_498 <= 1'h0;
    end else begin
      _T_498 <= _T_495;
    end
  end
endmodule
module FFType(
  input   clock,
  input   reset,
  input   io_in,
  input   io_init,
  output  io_out,
  input   io_enable
);
  wire  d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_10;
  wire  _GEN_0;
  wire  _GEN_1;
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? io_init : _T_10;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_10;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_10 = RetimeWrapper_io_out;
endmodule
module FF_2(
  input   clock,
  input   reset,
  input   io_in,
  input   io_init,
  output  io_out,
  input   io_enable
);
  wire  ff_clock;
  wire  ff_reset;
  wire  ff_io_in;
  wire  ff_io_init;
  wire  ff_io_out;
  wire  ff_io_enable;
  FFType ff (
    .clock(ff_clock),
    .reset(ff_reset),
    .io_in(ff_io_in),
    .io_init(ff_io_init),
    .io_out(ff_io_out),
    .io_enable(ff_io_enable)
  );
  assign io_out = ff_io_out;
  assign ff_io_in = io_in;
  assign ff_io_init = io_init;
  assign ff_io_enable = io_enable;
  assign ff_clock = clock;
  assign ff_reset = reset;
endmodule
module MuxVec(
  input  [63:0] io_ins_0_0_addr,
  input         io_ins_0_0_isWr,
  input  [15:0] io_ins_0_0_size,
  input  [63:0] io_ins_1_0_addr,
  input         io_ins_1_0_isWr,
  input  [15:0] io_ins_1_0_size,
  input         io_sel,
  output [63:0] io_out_0_addr,
  output        io_out_0_isWr,
  output [15:0] io_out_0_size
);
  wire [15:0] _GEN_0_0_size;
  wire [63:0] _GEN_4;
  wire  _GEN_5;
  wire [15:0] _GEN_7;
  wire  _GEN_2_0_isWr;
  wire [63:0] _GEN_3_0_addr;
  assign _GEN_4 = io_sel ? io_ins_1_0_addr : io_ins_0_0_addr;
  assign _GEN_5 = io_sel ? io_ins_1_0_isWr : io_ins_0_0_isWr;
  assign _GEN_7 = io_sel ? io_ins_1_0_size : io_ins_0_0_size;
  assign io_out_0_addr = _GEN_3_0_addr;
  assign io_out_0_isWr = _GEN_2_0_isWr;
  assign io_out_0_size = _GEN_0_0_size;
  assign _GEN_0_0_size = _GEN_7;
  assign _GEN_2_0_isWr = _GEN_5;
  assign _GEN_3_0_addr = _GEN_4;
endmodule
module FIFOArbiter(
  input         clock,
  input         reset,
  input  [63:0] io_fifo_0_deq_0_addr,
  input         io_fifo_0_deq_0_isWr,
  input  [15:0] io_fifo_0_deq_0_size,
  output        io_fifo_0_deqVld,
  input         io_fifo_0_empty,
  input         io_fifo_0_almostEmpty,
  input  [63:0] io_fifo_1_deq_0_addr,
  input         io_fifo_1_deq_0_isWr,
  input  [15:0] io_fifo_1_deq_0_size,
  output        io_fifo_1_deqVld,
  input         io_fifo_1_empty,
  output [63:0] io_deq_0_addr,
  output        io_deq_0_isWr,
  output [15:0] io_deq_0_size,
  input         io_deqVld,
  output        io_empty,
  output        io_tag
);
  wire  tagFF_clock;
  wire  tagFF_reset;
  wire  tagFF_io_in;
  wire  tagFF_io_init;
  wire  tagFF_io_out;
  wire  tagFF_io_enable;
  wire  tag;
  wire  _T_172;
  wire  _T_173;
  wire  _T_178;
  wire  _T_180;
  wire  _T_187;
  wire  _T_190;
  wire  _T_191;
  wire  _T_192;
  wire  _T_205_0;
  wire  _T_210_0;
  wire  _T_220;
  wire [63:0] MuxVec_io_ins_0_0_addr;
  wire  MuxVec_io_ins_0_0_isWr;
  wire [15:0] MuxVec_io_ins_0_0_size;
  wire [63:0] MuxVec_io_ins_1_0_addr;
  wire  MuxVec_io_ins_1_0_isWr;
  wire [15:0] MuxVec_io_ins_1_0_size;
  wire  MuxVec_io_sel;
  wire [63:0] MuxVec_io_out_0_addr;
  wire  MuxVec_io_out_0_isWr;
  wire [15:0] MuxVec_io_out_0_size;
  wire [63:0] _T_238_0_0_addr;
  wire  _T_238_0_0_isWr;
  wire [15:0] _T_238_0_0_size;
  wire [63:0] _T_238_1_0_addr;
  wire  _T_238_1_0_isWr;
  wire [15:0] _T_238_1_0_size;
  wire  _T_290;
  wire  _T_291;
  wire  _T_292;
  FF_2 tagFF (
    .clock(tagFF_clock),
    .reset(tagFF_reset),
    .io_in(tagFF_io_in),
    .io_init(tagFF_io_init),
    .io_out(tagFF_io_out),
    .io_enable(tagFF_io_enable)
  );
  MuxVec MuxVec (
    .io_ins_0_0_addr(MuxVec_io_ins_0_0_addr),
    .io_ins_0_0_isWr(MuxVec_io_ins_0_0_isWr),
    .io_ins_0_0_size(MuxVec_io_ins_0_0_size),
    .io_ins_1_0_addr(MuxVec_io_ins_1_0_addr),
    .io_ins_1_0_isWr(MuxVec_io_ins_1_0_isWr),
    .io_ins_1_0_size(MuxVec_io_ins_1_0_size),
    .io_sel(MuxVec_io_sel),
    .io_out_0_addr(MuxVec_io_out_0_addr),
    .io_out_0_isWr(MuxVec_io_out_0_isWr),
    .io_out_0_size(MuxVec_io_out_0_size)
  );
  assign tag = tagFF_io_out;
  assign _T_172 = tag == 1'h0;
  assign _T_173 = io_deqVld & _T_172;
  assign _T_178 = io_deqVld & tag;
  assign _T_180 = io_fifo_0_empty & io_fifo_1_empty;
  assign _T_187 = _T_172 & io_deqVld;
  assign _T_190 = _T_187 & io_fifo_0_almostEmpty;
  assign _T_191 = io_fifo_0_empty | _T_190;
  assign _T_192 = ~ _T_191;
  assign _T_210_0 = _T_180 ? 1'h0 : _T_205_0;
  assign _T_220 = _T_210_0 ? 1'h0 : 1'h1;
  assign _T_290 = tag ? io_fifo_1_empty : 1'h0;
  assign _T_291 = 1'h0 == tag;
  assign _T_292 = _T_291 ? io_fifo_0_empty : _T_290;
  assign io_fifo_0_deqVld = _T_173;
  assign io_fifo_1_deqVld = _T_178;
  assign io_deq_0_addr = MuxVec_io_out_0_addr;
  assign io_deq_0_isWr = MuxVec_io_out_0_isWr;
  assign io_deq_0_size = MuxVec_io_out_0_size;
  assign io_empty = _T_292;
  assign io_tag = tag;
  assign tagFF_io_in = _T_220;
  assign tagFF_io_init = 1'h0;
  assign tagFF_io_enable = io_deqVld;
  assign tagFF_clock = clock;
  assign tagFF_reset = reset;
  assign _T_205_0 = _T_192;
  assign MuxVec_io_ins_0_0_addr = _T_238_0_0_addr;
  assign MuxVec_io_ins_0_0_isWr = _T_238_0_0_isWr;
  assign MuxVec_io_ins_0_0_size = _T_238_0_0_size;
  assign MuxVec_io_ins_1_0_addr = _T_238_1_0_addr;
  assign MuxVec_io_ins_1_0_isWr = _T_238_1_0_isWr;
  assign MuxVec_io_ins_1_0_size = _T_238_1_0_size;
  assign MuxVec_io_sel = tag;
  assign _T_238_0_0_addr = io_fifo_0_deq_0_addr;
  assign _T_238_0_0_isWr = io_fifo_0_deq_0_isWr;
  assign _T_238_0_0_size = io_fifo_0_deq_0_size;
  assign _T_238_1_0_addr = io_fifo_1_deq_0_addr;
  assign _T_238_1_0_isWr = io_fifo_1_deq_0_isWr;
  assign _T_238_1_0_size = io_fifo_1_deq_0_size;
endmodule
module RetimeWrapper_7(
  input        clock,
  input        reset,
  input  [9:0] io_in,
  output [9:0] io_out
);
  wire [9:0] sr_out;
  wire [9:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(10), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FFType_1(
  input        clock,
  input        reset,
  input  [9:0] io_in,
  output [9:0] io_out,
  input        io_enable
);
  wire [9:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [9:0] RetimeWrapper_io_in;
  wire [9:0] RetimeWrapper_io_out;
  wire [9:0] _T_10;
  wire [9:0] _GEN_0;
  wire [9:0] _GEN_1;
  RetimeWrapper_7 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? 10'h0 : _T_10;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_10;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_10 = RetimeWrapper_io_out;
endmodule
module FF_3(
  input        clock,
  input        reset,
  input  [9:0] io_in,
  output [9:0] io_out,
  input        io_enable
);
  wire  ff_clock;
  wire  ff_reset;
  wire [9:0] ff_io_in;
  wire [9:0] ff_io_out;
  wire  ff_io_enable;
  FFType_1 ff (
    .clock(ff_clock),
    .reset(ff_reset),
    .io_in(ff_io_in),
    .io_out(ff_io_out),
    .io_enable(ff_io_enable)
  );
  assign io_out = ff_io_out;
  assign ff_io_in = io_in;
  assign ff_io_enable = io_enable;
  assign ff_clock = clock;
  assign ff_reset = reset;
endmodule
module UpDownCtr(
  input        clock,
  input        reset,
  input  [9:0] io_strideInc,
  input  [9:0] io_strideDec,
  input        io_inc,
  input        io_dec,
  output [9:0] io_out,
  output [9:0] io_nextInc,
  output [9:0] io_nextDec
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [9:0] reg$_io_in;
  wire [9:0] reg$_io_out;
  wire  reg$_io_enable;
  wire  _T_16;
  wire [9:0] incval;
  wire [9:0] decval;
  wire [10:0] _T_20;
  wire [10:0] _T_21;
  wire [9:0] incr;
  wire [10:0] _T_22;
  wire [9:0] newval;
  wire [10:0] _T_27;
  wire [9:0] _T_28;
  wire [10:0] _T_29;
  wire [10:0] _T_30;
  wire [9:0] _T_31;
  FF_3 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign _T_16 = io_inc | io_dec;
  assign incval = io_inc ? io_strideInc : 10'h0;
  assign decval = io_dec ? io_strideDec : 10'h0;
  assign _T_20 = incval - decval;
  assign _T_21 = $unsigned(_T_20);
  assign incr = _T_21[9:0];
  assign _T_22 = reg$_io_out + incr;
  assign newval = _T_22[9:0];
  assign _T_27 = reg$_io_out + io_strideInc;
  assign _T_28 = _T_27[9:0];
  assign _T_29 = reg$_io_out - io_strideDec;
  assign _T_30 = $unsigned(_T_29);
  assign _T_31 = _T_30[9:0];
  assign io_out = reg$_io_out;
  assign io_nextInc = _T_28;
  assign io_nextDec = _T_31;
  assign reg$_io_in = newval;
  assign reg$_io_enable = _T_16;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module Counter(
  input        clock,
  input        reset,
  input  [9:0] io_max,
  output [9:0] io_out,
  output [9:0] io_next,
  input        io_enable,
  output       io_done
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [9:0] reg$_io_in;
  wire [9:0] reg$_io_out;
  wire  reg$_io_enable;
  wire [10:0] count;
  wire [11:0] _T_12;
  wire [10:0] newval;
  wire [10:0] _GEN_1;
  wire  isMax;
  wire [10:0] next;
  wire  _T_14;
  FF_3 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out};
  assign _T_12 = count + 11'h1;
  assign newval = _T_12[10:0];
  assign _GEN_1 = {{1'd0}, io_max};
  assign isMax = newval >= _GEN_1;
  assign next = isMax ? 11'h0 : newval;
  assign _T_14 = io_enable & isMax;
  assign io_out = count[9:0];
  assign io_next = next[9:0];
  assign io_done = _T_14;
  assign reg$_io_in = next[9:0];
  assign reg$_io_enable = io_enable;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module Depulser(
  input   clock,
  input   reset,
  input   io_in,
  input   io_rst,
  output  io_out
);
  wire  r_clock;
  wire  r_reset;
  wire  r_io_in;
  wire  r_io_init;
  wire  r_io_out;
  wire  r_io_enable;
  wire  _T_6;
  wire  _T_8;
  FF_2 r (
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_init(r_io_init),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign _T_6 = io_rst ? 1'h0 : io_in;
  assign _T_8 = io_in | io_rst;
  assign io_out = r_io_out;
  assign r_io_in = _T_6;
  assign r_io_init = 1'h0;
  assign r_io_enable = _T_8;
  assign r_clock = clock;
  assign r_reset = reset;
endmodule
module CounterCore(
  input        clock,
  input        reset,
  output [9:0] io_out,
  output [9:0] io_next,
  input        io_enable,
  output       io_done,
  input  [9:0] io_config_max
);
  wire  counter_clock;
  wire  counter_reset;
  wire [9:0] counter_io_max;
  wire [9:0] counter_io_out;
  wire [9:0] counter_io_next;
  wire  counter_io_enable;
  wire  counter_io_done;
  wire  depulser_clock;
  wire  depulser_reset;
  wire  depulser_io_in;
  wire  depulser_io_rst;
  wire  depulser_io_out;
  Counter counter (
    .clock(counter_clock),
    .reset(counter_reset),
    .io_max(counter_io_max),
    .io_out(counter_io_out),
    .io_next(counter_io_next),
    .io_enable(counter_io_enable),
    .io_done(counter_io_done)
  );
  Depulser depulser (
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign io_out = counter_io_out;
  assign io_next = counter_io_next;
  assign io_done = counter_io_done;
  assign counter_io_max = io_config_max;
  assign counter_io_enable = io_enable;
  assign counter_clock = clock;
  assign counter_reset = reset;
  assign depulser_io_in = counter_io_done;
  assign depulser_io_rst = 1'h0;
  assign depulser_clock = clock;
  assign depulser_reset = reset;
endmodule
module CounterChainCore(
  input        clock,
  input        reset,
  output [9:0] io_out_1,
  output [9:0] io_next_1,
  input        io_enable_0,
  output       io_done_0
);
  wire  counters_0_clock;
  wire  counters_0_reset;
  wire [9:0] counters_0_io_out;
  wire [9:0] counters_0_io_next;
  wire  counters_0_io_enable;
  wire  counters_0_io_done;
  wire [9:0] counters_0_io_config_max;
  wire  counters_1_clock;
  wire  counters_1_reset;
  wire [9:0] counters_1_io_out;
  wire [9:0] counters_1_io_next;
  wire  counters_1_io_enable;
  wire  counters_1_io_done;
  wire [9:0] counters_1_io_config_max;
  wire  _T_69;
  CounterCore counters_0 (
    .clock(counters_0_clock),
    .reset(counters_0_reset),
    .io_out(counters_0_io_out),
    .io_next(counters_0_io_next),
    .io_enable(counters_0_io_enable),
    .io_done(counters_0_io_done),
    .io_config_max(counters_0_io_config_max)
  );
  CounterCore counters_1 (
    .clock(counters_1_clock),
    .reset(counters_1_reset),
    .io_out(counters_1_io_out),
    .io_next(counters_1_io_next),
    .io_enable(counters_1_io_enable),
    .io_done(counters_1_io_done),
    .io_config_max(counters_1_io_config_max)
  );
  assign _T_69 = counters_0_io_done;
  assign io_out_1 = counters_1_io_out;
  assign io_next_1 = counters_1_io_next;
  assign io_done_0 = counters_0_io_done;
  assign counters_0_io_enable = io_enable_0;
  assign counters_0_io_config_max = 10'h1;
  assign counters_0_clock = clock;
  assign counters_0_reset = reset;
  assign counters_1_io_enable = _T_69;
  assign counters_1_io_config_max = 10'h200;
  assign counters_1_clock = clock;
  assign counters_1_reset = reset;
endmodule
module SRAM(
  input         clock,
  input  [8:0]  io_raddr,
  input  [8:0]  io_waddr,
  output [63:0] io_rdata_addr,
  output        io_rdata_isWr,
  output [15:0] io_rdata_size
);
  wire [81:0] SRAMVerilogAWS_rdata;
  wire [81:0] SRAMVerilogAWS_wdata;
  wire  SRAMVerilogAWS_flow;
  wire  SRAMVerilogAWS_wen;
  wire  SRAMVerilogAWS_waddrEn;
  wire  SRAMVerilogAWS_raddrEn;
  wire [8:0] SRAMVerilogAWS_waddr;
  wire [8:0] SRAMVerilogAWS_raddr;
  wire  SRAMVerilogAWS_clk;
  wire [81:0] _T_22;
  wire [63:0] _T_24_addr;
  wire  _T_24_isWr;
  wire [15:0] _T_24_size;
  wire [81:0] _T_26;
  wire [15:0] _T_27;
  wire  _T_29;
  wire [63:0] _T_30;
  SRAMVerilogAWS #(.DWIDTH(82), .WORDS(512), .AWIDTH(9)) SRAMVerilogAWS (
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .flow(SRAMVerilogAWS_flow),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_22 = SRAMVerilogAWS_rdata;
  assign _T_27 = _T_26[15:0];
  assign _T_29 = _T_26[17];
  assign _T_30 = _T_26[81:18];
  assign io_rdata_addr = _T_24_addr;
  assign io_rdata_isWr = _T_24_isWr;
  assign io_rdata_size = _T_24_size;
  assign SRAMVerilogAWS_wdata = 82'h0;
  assign SRAMVerilogAWS_flow = 1'h1;
  assign SRAMVerilogAWS_wen = 1'h0;
  assign SRAMVerilogAWS_waddrEn = 1'h1;
  assign SRAMVerilogAWS_raddrEn = 1'h1;
  assign SRAMVerilogAWS_waddr = io_waddr;
  assign SRAMVerilogAWS_raddr = io_raddr;
  assign SRAMVerilogAWS_clk = clock;
  assign _T_24_addr = _T_30;
  assign _T_24_isWr = _T_29;
  assign _T_24_size = _T_27;
  assign _T_26 = _T_22;
endmodule
module MuxN_1(
  input  [63:0] io_ins_0_addr,
  input         io_ins_0_isWr,
  input  [15:0] io_ins_0_size,
  output [63:0] io_out_addr,
  output        io_out_isWr,
  output [15:0] io_out_size
);
  assign io_out_addr = io_ins_0_addr;
  assign io_out_isWr = io_ins_0_isWr;
  assign io_out_size = io_ins_0_size;
endmodule
module FIFOCore(
  input         clock,
  input         reset,
  output [63:0] io_deq_0_addr,
  output        io_deq_0_isWr,
  output [15:0] io_deq_0_size,
  input         io_deqVld,
  output        io_empty,
  output        io_almostEmpty
);
  wire  sizeUDC_clock;
  wire  sizeUDC_reset;
  wire [9:0] sizeUDC_io_strideInc;
  wire [9:0] sizeUDC_io_strideDec;
  wire  sizeUDC_io_inc;
  wire  sizeUDC_io_dec;
  wire [9:0] sizeUDC_io_out;
  wire [9:0] sizeUDC_io_nextInc;
  wire [9:0] sizeUDC_io_nextDec;
  wire  empty;
  wire  almostEmpty;
  wire  _T_35;
  wire  readEn;
  wire  wptr_clock;
  wire  wptr_reset;
  wire [9:0] wptr_io_out_1;
  wire [9:0] wptr_io_next_1;
  wire  wptr_io_enable_0;
  wire  wptr_io_done_0;
  wire  rptr_clock;
  wire  rptr_reset;
  wire [9:0] rptr_io_out_1;
  wire [9:0] rptr_io_next_1;
  wire  rptr_io_enable_0;
  wire  rptr_io_done_0;
  wire [9:0] nextHeadLocalAddr;
  wire  mems_0_0_clock;
  wire [8:0] mems_0_0_io_raddr;
  wire [8:0] mems_0_0_io_waddr;
  wire [63:0] mems_0_0_io_rdata_addr;
  wire  mems_0_0_io_rdata_isWr;
  wire [15:0] mems_0_0_io_rdata_size;
  wire [9:0] _T_79;
  wire [63:0] MuxN_io_ins_0_addr;
  wire  MuxN_io_ins_0_isWr;
  wire [15:0] MuxN_io_ins_0_size;
  wire [63:0] MuxN_io_out_addr;
  wire  MuxN_io_out_isWr;
  wire [15:0] MuxN_io_out_size;
  UpDownCtr sizeUDC (
    .clock(sizeUDC_clock),
    .reset(sizeUDC_reset),
    .io_strideInc(sizeUDC_io_strideInc),
    .io_strideDec(sizeUDC_io_strideDec),
    .io_inc(sizeUDC_io_inc),
    .io_dec(sizeUDC_io_dec),
    .io_out(sizeUDC_io_out),
    .io_nextInc(sizeUDC_io_nextInc),
    .io_nextDec(sizeUDC_io_nextDec)
  );
  CounterChainCore wptr (
    .clock(wptr_clock),
    .reset(wptr_reset),
    .io_out_1(wptr_io_out_1),
    .io_next_1(wptr_io_next_1),
    .io_enable_0(wptr_io_enable_0),
    .io_done_0(wptr_io_done_0)
  );
  CounterChainCore rptr (
    .clock(rptr_clock),
    .reset(rptr_reset),
    .io_out_1(rptr_io_out_1),
    .io_next_1(rptr_io_next_1),
    .io_enable_0(rptr_io_enable_0),
    .io_done_0(rptr_io_done_0)
  );
  SRAM mems_0_0 (
    .clock(mems_0_0_clock),
    .io_raddr(mems_0_0_io_raddr),
    .io_waddr(mems_0_0_io_waddr),
    .io_rdata_addr(mems_0_0_io_rdata_addr),
    .io_rdata_isWr(mems_0_0_io_rdata_isWr),
    .io_rdata_size(mems_0_0_io_rdata_size)
  );
  MuxN_1 MuxN (
    .io_ins_0_addr(MuxN_io_ins_0_addr),
    .io_ins_0_isWr(MuxN_io_ins_0_isWr),
    .io_ins_0_size(MuxN_io_ins_0_size),
    .io_out_addr(MuxN_io_out_addr),
    .io_out_isWr(MuxN_io_out_isWr),
    .io_out_size(MuxN_io_out_size)
  );
  assign empty = sizeUDC_io_out < 10'h1;
  assign almostEmpty = sizeUDC_io_nextDec < 10'h1;
  assign _T_35 = ~ empty;
  assign readEn = io_deqVld & _T_35;
  assign nextHeadLocalAddr = rptr_io_done_0 ? rptr_io_next_1 : rptr_io_out_1;
  assign _T_79 = readEn ? nextHeadLocalAddr : rptr_io_out_1;
  assign io_deq_0_addr = MuxN_io_out_addr;
  assign io_deq_0_isWr = MuxN_io_out_isWr;
  assign io_deq_0_size = MuxN_io_out_size;
  assign io_empty = empty;
  assign io_almostEmpty = almostEmpty;
  assign sizeUDC_io_strideInc = 10'h1;
  assign sizeUDC_io_strideDec = 10'h1;
  assign sizeUDC_io_inc = 1'h0;
  assign sizeUDC_io_dec = readEn;
  assign sizeUDC_clock = clock;
  assign sizeUDC_reset = reset;
  assign wptr_io_enable_0 = 1'h0;
  assign wptr_clock = clock;
  assign wptr_reset = reset;
  assign rptr_io_enable_0 = readEn;
  assign rptr_clock = clock;
  assign rptr_reset = reset;
  assign mems_0_0_io_raddr = _T_79[8:0];
  assign mems_0_0_io_waddr = wptr_io_out_1[8:0];
  assign mems_0_0_clock = clock;
  assign MuxN_io_ins_0_addr = mems_0_0_io_rdata_addr;
  assign MuxN_io_ins_0_isWr = mems_0_0_io_rdata_isWr;
  assign MuxN_io_ins_0_size = mems_0_0_io_rdata_size;
endmodule
module RetimeWrapper_25(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  output [31:0] io_out
);
  wire [31:0] sr_out;
  wire [31:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FFType_21(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  input  [31:0] io_init,
  output [31:0] io_out,
  input         io_enable
);
  wire [31:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [31:0] RetimeWrapper_io_in;
  wire [31:0] RetimeWrapper_io_out;
  wire [31:0] _T_10;
  wire [31:0] _GEN_0;
  wire [31:0] _GEN_1;
  RetimeWrapper_25 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? io_init : _T_10;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_10;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_10 = RetimeWrapper_io_out;
endmodule
module FF_23(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  input  [31:0] io_init,
  output [31:0] io_out,
  input         io_enable
);
  wire  ff_clock;
  wire  ff_reset;
  wire [31:0] ff_io_in;
  wire [31:0] ff_io_init;
  wire [31:0] ff_io_out;
  wire  ff_io_enable;
  FFType_21 ff (
    .clock(ff_clock),
    .reset(ff_reset),
    .io_in(ff_io_in),
    .io_init(ff_io_init),
    .io_out(ff_io_out),
    .io_enable(ff_io_enable)
  );
  assign io_out = ff_io_out;
  assign ff_io_in = io_in;
  assign ff_io_init = io_init;
  assign ff_io_enable = io_enable;
  assign ff_clock = clock;
  assign ff_reset = reset;
endmodule
module Counter_8(
  input         clock,
  input         reset,
  input  [31:0] io_max,
  output [31:0] io_out,
  input         io_enable,
  output        io_done
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [31:0] reg$_io_in;
  wire [31:0] reg$_io_init;
  wire [31:0] reg$_io_out;
  wire  reg$_io_enable;
  wire [32:0] count;
  wire [33:0] _T_12;
  wire [32:0] newval;
  wire [32:0] _GEN_1;
  wire  isMax;
  wire [32:0] next;
  wire  _T_14;
  FF_23 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_init(reg$_io_init),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out};
  assign _T_12 = count + 33'h1;
  assign newval = _T_12[32:0];
  assign _GEN_1 = {{1'd0}, io_max};
  assign isMax = newval >= _GEN_1;
  assign next = isMax ? 33'h0 : newval;
  assign _T_14 = io_enable & isMax;
  assign io_out = count[31:0];
  assign io_done = _T_14;
  assign reg$_io_in = next[31:0];
  assign reg$_io_init = 32'h0;
  assign reg$_io_enable = io_enable;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module MuxN_3(
  input   io_ins_0,
  output  io_out
);
  assign io_out = io_ins_0;
endmodule
module MuxN_4(
  input         io_ins_0_valid,
  input  [31:0] io_ins_0_bits_wdata_0,
  input  [31:0] io_ins_0_bits_wdata_1,
  input  [31:0] io_ins_0_bits_wdata_2,
  input  [31:0] io_ins_0_bits_wdata_3,
  input  [31:0] io_ins_0_bits_wdata_4,
  input  [31:0] io_ins_0_bits_wdata_5,
  input  [31:0] io_ins_0_bits_wdata_6,
  input  [31:0] io_ins_0_bits_wdata_7,
  input  [31:0] io_ins_0_bits_wdata_8,
  input  [31:0] io_ins_0_bits_wdata_9,
  input  [31:0] io_ins_0_bits_wdata_10,
  input  [31:0] io_ins_0_bits_wdata_11,
  input  [31:0] io_ins_0_bits_wdata_12,
  input  [31:0] io_ins_0_bits_wdata_13,
  input  [31:0] io_ins_0_bits_wdata_14,
  input  [31:0] io_ins_0_bits_wdata_15,
  input         io_ins_0_bits_wlast,
  output        io_out_valid,
  output [31:0] io_out_bits_wdata_0,
  output [31:0] io_out_bits_wdata_1,
  output [31:0] io_out_bits_wdata_2,
  output [31:0] io_out_bits_wdata_3,
  output [31:0] io_out_bits_wdata_4,
  output [31:0] io_out_bits_wdata_5,
  output [31:0] io_out_bits_wdata_6,
  output [31:0] io_out_bits_wdata_7,
  output [31:0] io_out_bits_wdata_8,
  output [31:0] io_out_bits_wdata_9,
  output [31:0] io_out_bits_wdata_10,
  output [31:0] io_out_bits_wdata_11,
  output [31:0] io_out_bits_wdata_12,
  output [31:0] io_out_bits_wdata_13,
  output [31:0] io_out_bits_wdata_14,
  output [31:0] io_out_bits_wdata_15,
  output        io_out_bits_wlast
);
  assign io_out_valid = io_ins_0_valid;
  assign io_out_bits_wdata_0 = io_ins_0_bits_wdata_0;
  assign io_out_bits_wdata_1 = io_ins_0_bits_wdata_1;
  assign io_out_bits_wdata_2 = io_ins_0_bits_wdata_2;
  assign io_out_bits_wdata_3 = io_ins_0_bits_wdata_3;
  assign io_out_bits_wdata_4 = io_ins_0_bits_wdata_4;
  assign io_out_bits_wdata_5 = io_ins_0_bits_wdata_5;
  assign io_out_bits_wdata_6 = io_ins_0_bits_wdata_6;
  assign io_out_bits_wdata_7 = io_ins_0_bits_wdata_7;
  assign io_out_bits_wdata_8 = io_ins_0_bits_wdata_8;
  assign io_out_bits_wdata_9 = io_ins_0_bits_wdata_9;
  assign io_out_bits_wdata_10 = io_ins_0_bits_wdata_10;
  assign io_out_bits_wdata_11 = io_ins_0_bits_wdata_11;
  assign io_out_bits_wdata_12 = io_ins_0_bits_wdata_12;
  assign io_out_bits_wdata_13 = io_ins_0_bits_wdata_13;
  assign io_out_bits_wdata_14 = io_ins_0_bits_wdata_14;
  assign io_out_bits_wdata_15 = io_ins_0_bits_wdata_15;
  assign io_out_bits_wlast = io_ins_0_bits_wlast;
endmodule
module MuxN_5(
  input   io_ins_0,
  input   io_ins_1,
  input   io_sel,
  output  io_out
);
  wire  _GEN_0;
  wire  _GEN_1;
  assign _GEN_1 = io_sel ? io_ins_1 : io_ins_0;
  assign io_out = _GEN_0;
  assign _GEN_0 = _GEN_1;
endmodule
module MuxN_6(
  input         io_ins_0_valid,
  input  [63:0] io_ins_0_bits_addr,
  input  [31:0] io_ins_0_bits_size,
  input         io_ins_0_bits_isWr,
  input  [25:0] io_ins_0_bits_tag_uid,
  input  [5:0]  io_ins_0_bits_tag_streamId,
  input         io_ins_1_valid,
  input  [63:0] io_ins_1_bits_addr,
  input  [31:0] io_ins_1_bits_size,
  input         io_ins_1_bits_isWr,
  input  [25:0] io_ins_1_bits_tag_uid,
  input  [5:0]  io_ins_1_bits_tag_streamId,
  input         io_sel,
  output        io_out_valid,
  output [63:0] io_out_bits_addr,
  output [31:0] io_out_bits_size,
  output        io_out_bits_isWr,
  output [25:0] io_out_bits_tag_uid,
  output [5:0]  io_out_bits_tag_streamId
);
  wire  _GEN_8;
  wire [63:0] _GEN_9;
  wire [31:0] _GEN_10;
  wire  _GEN_12;
  wire [25:0] _GEN_13;
  wire [5:0] _GEN_14;
  wire [5:0] _GEN_1_bits_tag_streamId;
  wire [25:0] _GEN_2_bits_tag_uid;
  wire  _GEN_3_bits_isWr;
  wire [31:0] _GEN_5_bits_size;
  wire [63:0] _GEN_6_bits_addr;
  wire  _GEN_7_valid;
  assign _GEN_8 = io_sel ? io_ins_1_valid : io_ins_0_valid;
  assign _GEN_9 = io_sel ? io_ins_1_bits_addr : io_ins_0_bits_addr;
  assign _GEN_10 = io_sel ? io_ins_1_bits_size : io_ins_0_bits_size;
  assign _GEN_12 = io_sel ? io_ins_1_bits_isWr : io_ins_0_bits_isWr;
  assign _GEN_13 = io_sel ? io_ins_1_bits_tag_uid : io_ins_0_bits_tag_uid;
  assign _GEN_14 = io_sel ? io_ins_1_bits_tag_streamId : io_ins_0_bits_tag_streamId;
  assign io_out_valid = _GEN_7_valid;
  assign io_out_bits_addr = _GEN_6_bits_addr;
  assign io_out_bits_size = _GEN_5_bits_size;
  assign io_out_bits_isWr = _GEN_3_bits_isWr;
  assign io_out_bits_tag_uid = _GEN_2_bits_tag_uid;
  assign io_out_bits_tag_streamId = _GEN_1_bits_tag_streamId;
  assign _GEN_1_bits_tag_streamId = _GEN_14;
  assign _GEN_2_bits_tag_uid = _GEN_13;
  assign _GEN_3_bits_isWr = _GEN_12;
  assign _GEN_5_bits_size = _GEN_10;
  assign _GEN_6_bits_addr = _GEN_9;
  assign _GEN_7_valid = _GEN_8;
endmodule
module RetimeWrapper_27(
  input        clock,
  input        reset,
  input  [5:0] io_in,
  output [5:0] io_out
);
  wire [5:0] sr_out;
  wire [5:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(6), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FFType_23(
  input        clock,
  input        reset,
  input  [5:0] io_in,
  input  [5:0] io_init,
  output [5:0] io_out,
  input        io_enable
);
  wire [5:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [5:0] RetimeWrapper_io_in;
  wire [5:0] RetimeWrapper_io_out;
  wire [5:0] _T_10;
  wire [5:0] _GEN_0;
  wire [5:0] _GEN_1;
  RetimeWrapper_27 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? io_init : _T_10;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_10;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_10 = RetimeWrapper_io_out;
endmodule
module FF_25(
  input        clock,
  input        reset,
  input  [5:0] io_in,
  input  [5:0] io_init,
  output [5:0] io_out,
  input        io_enable
);
  wire  ff_clock;
  wire  ff_reset;
  wire [5:0] ff_io_in;
  wire [5:0] ff_io_init;
  wire [5:0] ff_io_out;
  wire  ff_io_enable;
  FFType_23 ff (
    .clock(ff_clock),
    .reset(ff_reset),
    .io_in(ff_io_in),
    .io_init(ff_io_init),
    .io_out(ff_io_out),
    .io_enable(ff_io_enable)
  );
  assign io_out = ff_io_out;
  assign ff_io_in = io_in;
  assign ff_io_init = io_init;
  assign ff_io_enable = io_enable;
  assign ff_clock = clock;
  assign ff_reset = reset;
endmodule
module RetimeWrapper_28(
  input         clock,
  input         reset,
  input  [63:0] io_in,
  output [63:0] io_out
);
  wire [63:0] sr_out;
  wire [63:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FFType_24(
  input         clock,
  input         reset,
  input  [63:0] io_in,
  input  [63:0] io_init,
  output [63:0] io_out,
  input         io_enable
);
  wire [63:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [63:0] RetimeWrapper_io_in;
  wire [63:0] RetimeWrapper_io_out;
  wire [63:0] _T_10;
  wire [63:0] _GEN_0;
  wire [63:0] _GEN_1;
  RetimeWrapper_28 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? io_init : _T_10;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_10;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_10 = RetimeWrapper_io_out;
endmodule
module FF_26(
  input         clock,
  input         reset,
  input  [63:0] io_in,
  input  [63:0] io_init,
  output [63:0] io_out,
  input         io_enable
);
  wire  ff_clock;
  wire  ff_reset;
  wire [63:0] ff_io_in;
  wire [63:0] ff_io_init;
  wire [63:0] ff_io_out;
  wire  ff_io_enable;
  FFType_24 ff (
    .clock(ff_clock),
    .reset(ff_reset),
    .io_in(ff_io_in),
    .io_init(ff_io_init),
    .io_out(ff_io_out),
    .io_enable(ff_io_enable)
  );
  assign io_out = ff_io_out;
  assign ff_io_in = io_in;
  assign ff_io_init = io_init;
  assign ff_io_enable = io_enable;
  assign ff_clock = clock;
  assign ff_reset = reset;
endmodule
module RetimeWrapper_32(
  input         clock,
  input         reset,
  input  [15:0] io_in,
  output [15:0] io_out
);
  wire [15:0] sr_out;
  wire [15:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(16), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FFType_28(
  input         clock,
  input         reset,
  input  [15:0] io_in,
  output [15:0] io_out,
  input         io_enable
);
  wire [15:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [15:0] RetimeWrapper_io_in;
  wire [15:0] RetimeWrapper_io_out;
  wire [15:0] _T_10;
  wire [15:0] _GEN_0;
  wire [15:0] _GEN_1;
  RetimeWrapper_32 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? 16'hd6fd : _T_10;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_10;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_10 = RetimeWrapper_io_out;
endmodule
module FF_30(
  input         clock,
  input         reset,
  input  [15:0] io_in,
  output [15:0] io_out,
  input         io_enable
);
  wire  ff_clock;
  wire  ff_reset;
  wire [15:0] ff_io_in;
  wire [15:0] ff_io_out;
  wire  ff_io_enable;
  FFType_28 ff (
    .clock(ff_clock),
    .reset(ff_reset),
    .io_in(ff_io_in),
    .io_out(ff_io_out),
    .io_enable(ff_io_enable)
  );
  assign io_out = ff_io_out;
  assign ff_io_in = io_in;
  assign ff_io_enable = io_enable;
  assign ff_clock = clock;
  assign ff_reset = reset;
endmodule
module Counter_16(
  input        clock,
  input        reset,
  input  [5:0] io_max,
  output [5:0] io_out,
  output [5:0] io_next,
  input        io_enable,
  output       io_done
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [5:0] reg$_io_in;
  wire [5:0] reg$_io_init;
  wire [5:0] reg$_io_out;
  wire  reg$_io_enable;
  wire [6:0] count;
  wire [7:0] _T_12;
  wire [6:0] newval;
  wire [6:0] _GEN_1;
  wire  isMax;
  wire [6:0] next;
  wire  _T_14;
  FF_25 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_init(reg$_io_init),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out};
  assign _T_12 = count + 7'h1;
  assign newval = _T_12[6:0];
  assign _GEN_1 = {{1'd0}, io_max};
  assign isMax = newval >= _GEN_1;
  assign next = isMax ? 7'h0 : newval;
  assign _T_14 = io_enable & isMax;
  assign io_out = count[5:0];
  assign io_next = next[5:0];
  assign io_done = _T_14;
  assign reg$_io_in = next[5:0];
  assign reg$_io_init = 6'h0;
  assign reg$_io_enable = io_enable;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module CounterCore_8(
  input        clock,
  input        reset,
  output [5:0] io_out,
  output [5:0] io_next,
  input        io_enable,
  input  [5:0] io_config_max
);
  wire  counter_clock;
  wire  counter_reset;
  wire [5:0] counter_io_max;
  wire [5:0] counter_io_out;
  wire [5:0] counter_io_next;
  wire  counter_io_enable;
  wire  counter_io_done;
  wire  depulser_clock;
  wire  depulser_reset;
  wire  depulser_io_in;
  wire  depulser_io_rst;
  wire  depulser_io_out;
  Counter_16 counter (
    .clock(counter_clock),
    .reset(counter_reset),
    .io_max(counter_io_max),
    .io_out(counter_io_out),
    .io_next(counter_io_next),
    .io_enable(counter_io_enable),
    .io_done(counter_io_done)
  );
  Depulser depulser (
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign io_out = counter_io_out;
  assign io_next = counter_io_next;
  assign counter_io_max = io_config_max;
  assign counter_io_enable = io_enable;
  assign counter_clock = clock;
  assign counter_reset = reset;
  assign depulser_io_in = counter_io_done;
  assign depulser_io_rst = 1'h0;
  assign depulser_clock = clock;
  assign depulser_reset = reset;
endmodule
module CounterChainCore_4(
  input        clock,
  input        reset,
  output [5:0] io_out_0,
  output [5:0] io_out_1,
  output [5:0] io_next_0,
  output [5:0] io_next_1,
  input        io_enable_1
);
  wire  counters_0_clock;
  wire  counters_0_reset;
  wire [5:0] counters_0_io_out;
  wire [5:0] counters_0_io_next;
  wire  counters_0_io_enable;
  wire [5:0] counters_0_io_config_max;
  wire  counters_1_clock;
  wire  counters_1_reset;
  wire [5:0] counters_1_io_out;
  wire [5:0] counters_1_io_next;
  wire  counters_1_io_enable;
  wire [5:0] counters_1_io_config_max;
  CounterCore_8 counters_0 (
    .clock(counters_0_clock),
    .reset(counters_0_reset),
    .io_out(counters_0_io_out),
    .io_next(counters_0_io_next),
    .io_enable(counters_0_io_enable),
    .io_config_max(counters_0_io_config_max)
  );
  CounterCore_8 counters_1 (
    .clock(counters_1_clock),
    .reset(counters_1_reset),
    .io_out(counters_1_io_out),
    .io_next(counters_1_io_next),
    .io_enable(counters_1_io_enable),
    .io_config_max(counters_1_io_config_max)
  );
  assign io_out_0 = counters_0_io_out;
  assign io_out_1 = counters_1_io_out;
  assign io_next_0 = counters_0_io_next;
  assign io_next_1 = counters_1_io_next;
  assign counters_0_io_enable = 1'h0;
  assign counters_0_io_config_max = 6'h10;
  assign counters_0_clock = clock;
  assign counters_0_reset = reset;
  assign counters_1_io_enable = io_enable_1;
  assign counters_1_io_config_max = 6'h20;
  assign counters_1_clock = clock;
  assign counters_1_reset = reset;
endmodule
module SRAM_2(
  input         clock,
  input         reset,
  input  [4:0]  io_raddr,
  input         io_wen,
  input  [4:0]  io_waddr,
  input  [31:0] io_wdata,
  output [31:0] io_rdata
);
  wire [31:0] SRAMVerilogAWS_rdata;
  wire [31:0] SRAMVerilogAWS_wdata;
  wire  SRAMVerilogAWS_flow;
  wire  SRAMVerilogAWS_wen;
  wire  SRAMVerilogAWS_waddrEn;
  wire  SRAMVerilogAWS_raddrEn;
  wire [4:0] SRAMVerilogAWS_waddr;
  wire [4:0] SRAMVerilogAWS_raddr;
  wire  SRAMVerilogAWS_clk;
  wire  _T_8;
  wire  _T_9;
  reg  _T_12;
  reg [31:0] _RAND_0;
  reg [31:0] _T_15;
  reg [31:0] _RAND_1;
  wire [31:0] _T_16;
  wire [31:0] _T_18;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(32), .AWIDTH(5)) SRAMVerilogAWS (
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .flow(SRAMVerilogAWS_flow),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_8 = io_raddr == io_waddr;
  assign _T_9 = io_wen & _T_8;
  assign _T_16 = _T_12 ? _T_15 : SRAMVerilogAWS_rdata;
  assign io_rdata = _T_18;
  assign SRAMVerilogAWS_wdata = io_wdata;
  assign SRAMVerilogAWS_flow = 1'h1;
  assign SRAMVerilogAWS_wen = io_wen;
  assign SRAMVerilogAWS_waddrEn = 1'h1;
  assign SRAMVerilogAWS_raddrEn = 1'h1;
  assign SRAMVerilogAWS_waddr = io_waddr;
  assign SRAMVerilogAWS_raddr = io_raddr;
  assign SRAMVerilogAWS_clk = clock;
  assign _T_18 = _T_16;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_12 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_15 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_12 <= 1'h0;
    end else begin
      _T_12 <= _T_9;
    end
    if (reset) begin
      _T_15 <= 32'h0;
    end else begin
      _T_15 <= io_wdata;
    end
  end
endmodule
module MuxN_14(
  input  [31:0] io_ins_0,
  output [31:0] io_out
);
  wire [31:0] _GEN_0;
  assign io_out = _GEN_0;
  assign _GEN_0 = io_ins_0;
endmodule
module RetimeWrapper_48(
  input        clock,
  input        reset,
  input  [3:0] io_in
);
  wire [3:0] sr_out;
  wire [3:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(4), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FFType_44(
  input        clock,
  input        reset,
  input  [3:0] io_in
);
  wire [3:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [3:0] RetimeWrapper_io_in;
  RetimeWrapper_48 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in)
  );
  assign d = io_in;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
endmodule
module FF_46(
  input        clock,
  input        reset,
  input  [3:0] io_in
);
  wire  ff_clock;
  wire  ff_reset;
  wire [3:0] ff_io_in;
  FFType_44 ff (
    .clock(ff_clock),
    .reset(ff_reset),
    .io_in(ff_io_in)
  );
  assign ff_io_in = io_in;
  assign ff_clock = clock;
  assign ff_reset = reset;
endmodule
module FIFOCore_2(
  input         clock,
  input         reset,
  input  [31:0] io_enq_0,
  input  [31:0] io_enq_1,
  input  [31:0] io_enq_2,
  input  [31:0] io_enq_3,
  input  [31:0] io_enq_4,
  input  [31:0] io_enq_5,
  input  [31:0] io_enq_6,
  input  [31:0] io_enq_7,
  input  [31:0] io_enq_8,
  input  [31:0] io_enq_9,
  input  [31:0] io_enq_10,
  input  [31:0] io_enq_11,
  input  [31:0] io_enq_12,
  input  [31:0] io_enq_13,
  input  [31:0] io_enq_14,
  input  [31:0] io_enq_15,
  input         io_enqVld,
  output [31:0] io_deq_0,
  output [31:0] io_deq_1,
  output [31:0] io_deq_2,
  output [31:0] io_deq_3,
  output [31:0] io_deq_4,
  output [31:0] io_deq_5,
  output [31:0] io_deq_6,
  output [31:0] io_deq_7,
  output [31:0] io_deq_8,
  output [31:0] io_deq_9,
  output [31:0] io_deq_10,
  output [31:0] io_deq_11,
  output [31:0] io_deq_12,
  output [31:0] io_deq_13,
  output [31:0] io_deq_14,
  output [31:0] io_deq_15,
  input         io_deqVld,
  output        io_full,
  output        io_empty,
  output        io_almostFull,
  output        io_almostEmpty
);
  wire  sizeUDC_clock;
  wire  sizeUDC_reset;
  wire [9:0] sizeUDC_io_strideInc;
  wire [9:0] sizeUDC_io_strideDec;
  wire  sizeUDC_io_inc;
  wire  sizeUDC_io_dec;
  wire [9:0] sizeUDC_io_out;
  wire [9:0] sizeUDC_io_nextInc;
  wire [9:0] sizeUDC_io_nextDec;
  wire [10:0] _T_51;
  wire [10:0] _T_52;
  wire [9:0] remainingSlots;
  wire [10:0] _T_54;
  wire [10:0] _T_55;
  wire [9:0] nextRemainingSlots;
  wire  empty;
  wire  almostEmpty;
  wire  full;
  wire  almostFull;
  wire  _T_64;
  wire  writeEn;
  wire  _T_65;
  wire  readEn;
  wire  wptr_clock;
  wire  wptr_reset;
  wire [5:0] wptr_io_out_0;
  wire [5:0] wptr_io_out_1;
  wire [5:0] wptr_io_next_0;
  wire [5:0] wptr_io_next_1;
  wire  wptr_io_enable_1;
  wire  rptr_clock;
  wire  rptr_reset;
  wire [5:0] rptr_io_out_0;
  wire [5:0] rptr_io_out_1;
  wire [5:0] rptr_io_next_0;
  wire [5:0] rptr_io_next_1;
  wire  rptr_io_enable_1;
  wire [5:0] nextHeadLocalAddr;
  wire  mems_0_0_clock;
  wire  mems_0_0_reset;
  wire [4:0] mems_0_0_io_raddr;
  wire  mems_0_0_io_wen;
  wire [4:0] mems_0_0_io_waddr;
  wire [31:0] mems_0_0_io_wdata;
  wire [31:0] mems_0_0_io_rdata;
  wire  mems_0_1_clock;
  wire  mems_0_1_reset;
  wire [4:0] mems_0_1_io_raddr;
  wire  mems_0_1_io_wen;
  wire [4:0] mems_0_1_io_waddr;
  wire [31:0] mems_0_1_io_wdata;
  wire [31:0] mems_0_1_io_rdata;
  wire  mems_0_2_clock;
  wire  mems_0_2_reset;
  wire [4:0] mems_0_2_io_raddr;
  wire  mems_0_2_io_wen;
  wire [4:0] mems_0_2_io_waddr;
  wire [31:0] mems_0_2_io_wdata;
  wire [31:0] mems_0_2_io_rdata;
  wire  mems_0_3_clock;
  wire  mems_0_3_reset;
  wire [4:0] mems_0_3_io_raddr;
  wire  mems_0_3_io_wen;
  wire [4:0] mems_0_3_io_waddr;
  wire [31:0] mems_0_3_io_wdata;
  wire [31:0] mems_0_3_io_rdata;
  wire  mems_0_4_clock;
  wire  mems_0_4_reset;
  wire [4:0] mems_0_4_io_raddr;
  wire  mems_0_4_io_wen;
  wire [4:0] mems_0_4_io_waddr;
  wire [31:0] mems_0_4_io_wdata;
  wire [31:0] mems_0_4_io_rdata;
  wire  mems_0_5_clock;
  wire  mems_0_5_reset;
  wire [4:0] mems_0_5_io_raddr;
  wire  mems_0_5_io_wen;
  wire [4:0] mems_0_5_io_waddr;
  wire [31:0] mems_0_5_io_wdata;
  wire [31:0] mems_0_5_io_rdata;
  wire  mems_0_6_clock;
  wire  mems_0_6_reset;
  wire [4:0] mems_0_6_io_raddr;
  wire  mems_0_6_io_wen;
  wire [4:0] mems_0_6_io_waddr;
  wire [31:0] mems_0_6_io_wdata;
  wire [31:0] mems_0_6_io_rdata;
  wire  mems_0_7_clock;
  wire  mems_0_7_reset;
  wire [4:0] mems_0_7_io_raddr;
  wire  mems_0_7_io_wen;
  wire [4:0] mems_0_7_io_waddr;
  wire [31:0] mems_0_7_io_wdata;
  wire [31:0] mems_0_7_io_rdata;
  wire  mems_0_8_clock;
  wire  mems_0_8_reset;
  wire [4:0] mems_0_8_io_raddr;
  wire  mems_0_8_io_wen;
  wire [4:0] mems_0_8_io_waddr;
  wire [31:0] mems_0_8_io_wdata;
  wire [31:0] mems_0_8_io_rdata;
  wire  mems_0_9_clock;
  wire  mems_0_9_reset;
  wire [4:0] mems_0_9_io_raddr;
  wire  mems_0_9_io_wen;
  wire [4:0] mems_0_9_io_waddr;
  wire [31:0] mems_0_9_io_wdata;
  wire [31:0] mems_0_9_io_rdata;
  wire  mems_0_10_clock;
  wire  mems_0_10_reset;
  wire [4:0] mems_0_10_io_raddr;
  wire  mems_0_10_io_wen;
  wire [4:0] mems_0_10_io_waddr;
  wire [31:0] mems_0_10_io_wdata;
  wire [31:0] mems_0_10_io_rdata;
  wire  mems_0_11_clock;
  wire  mems_0_11_reset;
  wire [4:0] mems_0_11_io_raddr;
  wire  mems_0_11_io_wen;
  wire [4:0] mems_0_11_io_waddr;
  wire [31:0] mems_0_11_io_wdata;
  wire [31:0] mems_0_11_io_rdata;
  wire  mems_0_12_clock;
  wire  mems_0_12_reset;
  wire [4:0] mems_0_12_io_raddr;
  wire  mems_0_12_io_wen;
  wire [4:0] mems_0_12_io_waddr;
  wire [31:0] mems_0_12_io_wdata;
  wire [31:0] mems_0_12_io_rdata;
  wire  mems_0_13_clock;
  wire  mems_0_13_reset;
  wire [4:0] mems_0_13_io_raddr;
  wire  mems_0_13_io_wen;
  wire [4:0] mems_0_13_io_waddr;
  wire [31:0] mems_0_13_io_wdata;
  wire [31:0] mems_0_13_io_rdata;
  wire  mems_0_14_clock;
  wire  mems_0_14_reset;
  wire [4:0] mems_0_14_io_raddr;
  wire  mems_0_14_io_wen;
  wire [4:0] mems_0_14_io_waddr;
  wire [31:0] mems_0_14_io_wdata;
  wire [31:0] mems_0_14_io_rdata;
  wire  mems_0_15_clock;
  wire  mems_0_15_reset;
  wire [4:0] mems_0_15_io_raddr;
  wire  mems_0_15_io_wen;
  wire [4:0] mems_0_15_io_waddr;
  wire [31:0] mems_0_15_io_wdata;
  wire [31:0] mems_0_15_io_rdata;
  wire [31:0] wdata_0;
  wire [31:0] wdata_1;
  wire [31:0] wdata_2;
  wire [31:0] wdata_3;
  wire [31:0] wdata_4;
  wire [31:0] wdata_5;
  wire [31:0] wdata_6;
  wire [31:0] wdata_7;
  wire [31:0] wdata_8;
  wire [31:0] wdata_9;
  wire [31:0] wdata_10;
  wire [31:0] wdata_11;
  wire [31:0] wdata_12;
  wire [31:0] wdata_13;
  wire [31:0] wdata_14;
  wire [31:0] wdata_15;
  wire [5:0] _T_154;
  wire [31:0] MuxN_io_ins_0;
  wire [31:0] MuxN_io_out;
  wire  FF_clock;
  wire  FF_reset;
  wire [3:0] FF_io_in;
  wire [5:0] _T_159;
  UpDownCtr sizeUDC (
    .clock(sizeUDC_clock),
    .reset(sizeUDC_reset),
    .io_strideInc(sizeUDC_io_strideInc),
    .io_strideDec(sizeUDC_io_strideDec),
    .io_inc(sizeUDC_io_inc),
    .io_dec(sizeUDC_io_dec),
    .io_out(sizeUDC_io_out),
    .io_nextInc(sizeUDC_io_nextInc),
    .io_nextDec(sizeUDC_io_nextDec)
  );
  CounterChainCore_4 wptr (
    .clock(wptr_clock),
    .reset(wptr_reset),
    .io_out_0(wptr_io_out_0),
    .io_out_1(wptr_io_out_1),
    .io_next_0(wptr_io_next_0),
    .io_next_1(wptr_io_next_1),
    .io_enable_1(wptr_io_enable_1)
  );
  CounterChainCore_4 rptr (
    .clock(rptr_clock),
    .reset(rptr_reset),
    .io_out_0(rptr_io_out_0),
    .io_out_1(rptr_io_out_1),
    .io_next_0(rptr_io_next_0),
    .io_next_1(rptr_io_next_1),
    .io_enable_1(rptr_io_enable_1)
  );
  SRAM_2 mems_0_0 (
    .clock(mems_0_0_clock),
    .reset(mems_0_0_reset),
    .io_raddr(mems_0_0_io_raddr),
    .io_wen(mems_0_0_io_wen),
    .io_waddr(mems_0_0_io_waddr),
    .io_wdata(mems_0_0_io_wdata),
    .io_rdata(mems_0_0_io_rdata)
  );
  SRAM_2 mems_0_1 (
    .clock(mems_0_1_clock),
    .reset(mems_0_1_reset),
    .io_raddr(mems_0_1_io_raddr),
    .io_wen(mems_0_1_io_wen),
    .io_waddr(mems_0_1_io_waddr),
    .io_wdata(mems_0_1_io_wdata),
    .io_rdata(mems_0_1_io_rdata)
  );
  SRAM_2 mems_0_2 (
    .clock(mems_0_2_clock),
    .reset(mems_0_2_reset),
    .io_raddr(mems_0_2_io_raddr),
    .io_wen(mems_0_2_io_wen),
    .io_waddr(mems_0_2_io_waddr),
    .io_wdata(mems_0_2_io_wdata),
    .io_rdata(mems_0_2_io_rdata)
  );
  SRAM_2 mems_0_3 (
    .clock(mems_0_3_clock),
    .reset(mems_0_3_reset),
    .io_raddr(mems_0_3_io_raddr),
    .io_wen(mems_0_3_io_wen),
    .io_waddr(mems_0_3_io_waddr),
    .io_wdata(mems_0_3_io_wdata),
    .io_rdata(mems_0_3_io_rdata)
  );
  SRAM_2 mems_0_4 (
    .clock(mems_0_4_clock),
    .reset(mems_0_4_reset),
    .io_raddr(mems_0_4_io_raddr),
    .io_wen(mems_0_4_io_wen),
    .io_waddr(mems_0_4_io_waddr),
    .io_wdata(mems_0_4_io_wdata),
    .io_rdata(mems_0_4_io_rdata)
  );
  SRAM_2 mems_0_5 (
    .clock(mems_0_5_clock),
    .reset(mems_0_5_reset),
    .io_raddr(mems_0_5_io_raddr),
    .io_wen(mems_0_5_io_wen),
    .io_waddr(mems_0_5_io_waddr),
    .io_wdata(mems_0_5_io_wdata),
    .io_rdata(mems_0_5_io_rdata)
  );
  SRAM_2 mems_0_6 (
    .clock(mems_0_6_clock),
    .reset(mems_0_6_reset),
    .io_raddr(mems_0_6_io_raddr),
    .io_wen(mems_0_6_io_wen),
    .io_waddr(mems_0_6_io_waddr),
    .io_wdata(mems_0_6_io_wdata),
    .io_rdata(mems_0_6_io_rdata)
  );
  SRAM_2 mems_0_7 (
    .clock(mems_0_7_clock),
    .reset(mems_0_7_reset),
    .io_raddr(mems_0_7_io_raddr),
    .io_wen(mems_0_7_io_wen),
    .io_waddr(mems_0_7_io_waddr),
    .io_wdata(mems_0_7_io_wdata),
    .io_rdata(mems_0_7_io_rdata)
  );
  SRAM_2 mems_0_8 (
    .clock(mems_0_8_clock),
    .reset(mems_0_8_reset),
    .io_raddr(mems_0_8_io_raddr),
    .io_wen(mems_0_8_io_wen),
    .io_waddr(mems_0_8_io_waddr),
    .io_wdata(mems_0_8_io_wdata),
    .io_rdata(mems_0_8_io_rdata)
  );
  SRAM_2 mems_0_9 (
    .clock(mems_0_9_clock),
    .reset(mems_0_9_reset),
    .io_raddr(mems_0_9_io_raddr),
    .io_wen(mems_0_9_io_wen),
    .io_waddr(mems_0_9_io_waddr),
    .io_wdata(mems_0_9_io_wdata),
    .io_rdata(mems_0_9_io_rdata)
  );
  SRAM_2 mems_0_10 (
    .clock(mems_0_10_clock),
    .reset(mems_0_10_reset),
    .io_raddr(mems_0_10_io_raddr),
    .io_wen(mems_0_10_io_wen),
    .io_waddr(mems_0_10_io_waddr),
    .io_wdata(mems_0_10_io_wdata),
    .io_rdata(mems_0_10_io_rdata)
  );
  SRAM_2 mems_0_11 (
    .clock(mems_0_11_clock),
    .reset(mems_0_11_reset),
    .io_raddr(mems_0_11_io_raddr),
    .io_wen(mems_0_11_io_wen),
    .io_waddr(mems_0_11_io_waddr),
    .io_wdata(mems_0_11_io_wdata),
    .io_rdata(mems_0_11_io_rdata)
  );
  SRAM_2 mems_0_12 (
    .clock(mems_0_12_clock),
    .reset(mems_0_12_reset),
    .io_raddr(mems_0_12_io_raddr),
    .io_wen(mems_0_12_io_wen),
    .io_waddr(mems_0_12_io_waddr),
    .io_wdata(mems_0_12_io_wdata),
    .io_rdata(mems_0_12_io_rdata)
  );
  SRAM_2 mems_0_13 (
    .clock(mems_0_13_clock),
    .reset(mems_0_13_reset),
    .io_raddr(mems_0_13_io_raddr),
    .io_wen(mems_0_13_io_wen),
    .io_waddr(mems_0_13_io_waddr),
    .io_wdata(mems_0_13_io_wdata),
    .io_rdata(mems_0_13_io_rdata)
  );
  SRAM_2 mems_0_14 (
    .clock(mems_0_14_clock),
    .reset(mems_0_14_reset),
    .io_raddr(mems_0_14_io_raddr),
    .io_wen(mems_0_14_io_wen),
    .io_waddr(mems_0_14_io_waddr),
    .io_wdata(mems_0_14_io_wdata),
    .io_rdata(mems_0_14_io_rdata)
  );
  SRAM_2 mems_0_15 (
    .clock(mems_0_15_clock),
    .reset(mems_0_15_reset),
    .io_raddr(mems_0_15_io_raddr),
    .io_wen(mems_0_15_io_wen),
    .io_waddr(mems_0_15_io_waddr),
    .io_wdata(mems_0_15_io_wdata),
    .io_rdata(mems_0_15_io_rdata)
  );
  MuxN_14 MuxN (
    .io_ins_0(MuxN_io_ins_0),
    .io_out(MuxN_io_out)
  );
  FF_46 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_in(FF_io_in)
  );
  assign _T_51 = 10'h200 - sizeUDC_io_out;
  assign _T_52 = $unsigned(_T_51);
  assign remainingSlots = _T_52[9:0];
  assign _T_54 = 10'h200 - sizeUDC_io_nextInc;
  assign _T_55 = $unsigned(_T_54);
  assign nextRemainingSlots = _T_55[9:0];
  assign empty = sizeUDC_io_out < 10'h10;
  assign almostEmpty = sizeUDC_io_nextDec < 10'h10;
  assign full = remainingSlots < 10'h10;
  assign almostFull = nextRemainingSlots < 10'h10;
  assign _T_64 = ~ full;
  assign writeEn = io_enqVld & _T_64;
  assign _T_65 = ~ empty;
  assign readEn = io_deqVld & _T_65;
  assign nextHeadLocalAddr = rptr_io_next_1;
  assign _T_154 = readEn ? nextHeadLocalAddr : rptr_io_out_1;
  assign _T_159 = readEn ? rptr_io_next_0 : rptr_io_out_0;
  assign io_deq_0 = MuxN_io_out;
  assign io_deq_1 = mems_0_1_io_rdata;
  assign io_deq_2 = mems_0_2_io_rdata;
  assign io_deq_3 = mems_0_3_io_rdata;
  assign io_deq_4 = mems_0_4_io_rdata;
  assign io_deq_5 = mems_0_5_io_rdata;
  assign io_deq_6 = mems_0_6_io_rdata;
  assign io_deq_7 = mems_0_7_io_rdata;
  assign io_deq_8 = mems_0_8_io_rdata;
  assign io_deq_9 = mems_0_9_io_rdata;
  assign io_deq_10 = mems_0_10_io_rdata;
  assign io_deq_11 = mems_0_11_io_rdata;
  assign io_deq_12 = mems_0_12_io_rdata;
  assign io_deq_13 = mems_0_13_io_rdata;
  assign io_deq_14 = mems_0_14_io_rdata;
  assign io_deq_15 = mems_0_15_io_rdata;
  assign io_full = full;
  assign io_empty = empty;
  assign io_almostFull = almostFull;
  assign io_almostEmpty = almostEmpty;
  assign sizeUDC_io_strideInc = 10'h10;
  assign sizeUDC_io_strideDec = 10'h10;
  assign sizeUDC_io_inc = writeEn;
  assign sizeUDC_io_dec = readEn;
  assign sizeUDC_clock = clock;
  assign sizeUDC_reset = reset;
  assign wptr_io_enable_1 = writeEn;
  assign wptr_clock = clock;
  assign wptr_reset = reset;
  assign rptr_io_enable_1 = readEn;
  assign rptr_clock = clock;
  assign rptr_reset = reset;
  assign mems_0_0_io_raddr = _T_154[4:0];
  assign mems_0_0_io_wen = writeEn;
  assign mems_0_0_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_0_io_wdata = wdata_0;
  assign mems_0_0_clock = clock;
  assign mems_0_0_reset = reset;
  assign mems_0_1_io_raddr = _T_154[4:0];
  assign mems_0_1_io_wen = writeEn;
  assign mems_0_1_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_1_io_wdata = wdata_1;
  assign mems_0_1_clock = clock;
  assign mems_0_1_reset = reset;
  assign mems_0_2_io_raddr = _T_154[4:0];
  assign mems_0_2_io_wen = writeEn;
  assign mems_0_2_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_2_io_wdata = wdata_2;
  assign mems_0_2_clock = clock;
  assign mems_0_2_reset = reset;
  assign mems_0_3_io_raddr = _T_154[4:0];
  assign mems_0_3_io_wen = writeEn;
  assign mems_0_3_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_3_io_wdata = wdata_3;
  assign mems_0_3_clock = clock;
  assign mems_0_3_reset = reset;
  assign mems_0_4_io_raddr = _T_154[4:0];
  assign mems_0_4_io_wen = writeEn;
  assign mems_0_4_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_4_io_wdata = wdata_4;
  assign mems_0_4_clock = clock;
  assign mems_0_4_reset = reset;
  assign mems_0_5_io_raddr = _T_154[4:0];
  assign mems_0_5_io_wen = writeEn;
  assign mems_0_5_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_5_io_wdata = wdata_5;
  assign mems_0_5_clock = clock;
  assign mems_0_5_reset = reset;
  assign mems_0_6_io_raddr = _T_154[4:0];
  assign mems_0_6_io_wen = writeEn;
  assign mems_0_6_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_6_io_wdata = wdata_6;
  assign mems_0_6_clock = clock;
  assign mems_0_6_reset = reset;
  assign mems_0_7_io_raddr = _T_154[4:0];
  assign mems_0_7_io_wen = writeEn;
  assign mems_0_7_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_7_io_wdata = wdata_7;
  assign mems_0_7_clock = clock;
  assign mems_0_7_reset = reset;
  assign mems_0_8_io_raddr = _T_154[4:0];
  assign mems_0_8_io_wen = writeEn;
  assign mems_0_8_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_8_io_wdata = wdata_8;
  assign mems_0_8_clock = clock;
  assign mems_0_8_reset = reset;
  assign mems_0_9_io_raddr = _T_154[4:0];
  assign mems_0_9_io_wen = writeEn;
  assign mems_0_9_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_9_io_wdata = wdata_9;
  assign mems_0_9_clock = clock;
  assign mems_0_9_reset = reset;
  assign mems_0_10_io_raddr = _T_154[4:0];
  assign mems_0_10_io_wen = writeEn;
  assign mems_0_10_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_10_io_wdata = wdata_10;
  assign mems_0_10_clock = clock;
  assign mems_0_10_reset = reset;
  assign mems_0_11_io_raddr = _T_154[4:0];
  assign mems_0_11_io_wen = writeEn;
  assign mems_0_11_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_11_io_wdata = wdata_11;
  assign mems_0_11_clock = clock;
  assign mems_0_11_reset = reset;
  assign mems_0_12_io_raddr = _T_154[4:0];
  assign mems_0_12_io_wen = writeEn;
  assign mems_0_12_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_12_io_wdata = wdata_12;
  assign mems_0_12_clock = clock;
  assign mems_0_12_reset = reset;
  assign mems_0_13_io_raddr = _T_154[4:0];
  assign mems_0_13_io_wen = writeEn;
  assign mems_0_13_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_13_io_wdata = wdata_13;
  assign mems_0_13_clock = clock;
  assign mems_0_13_reset = reset;
  assign mems_0_14_io_raddr = _T_154[4:0];
  assign mems_0_14_io_wen = writeEn;
  assign mems_0_14_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_14_io_wdata = wdata_14;
  assign mems_0_14_clock = clock;
  assign mems_0_14_reset = reset;
  assign mems_0_15_io_raddr = _T_154[4:0];
  assign mems_0_15_io_wen = writeEn;
  assign mems_0_15_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_15_io_wdata = wdata_15;
  assign mems_0_15_clock = clock;
  assign mems_0_15_reset = reset;
  assign wdata_0 = io_enq_0;
  assign wdata_1 = io_enq_1;
  assign wdata_2 = io_enq_2;
  assign wdata_3 = io_enq_3;
  assign wdata_4 = io_enq_4;
  assign wdata_5 = io_enq_5;
  assign wdata_6 = io_enq_6;
  assign wdata_7 = io_enq_7;
  assign wdata_8 = io_enq_8;
  assign wdata_9 = io_enq_9;
  assign wdata_10 = io_enq_10;
  assign wdata_11 = io_enq_11;
  assign wdata_12 = io_enq_12;
  assign wdata_13 = io_enq_13;
  assign wdata_14 = io_enq_14;
  assign wdata_15 = io_enq_15;
  assign MuxN_io_ins_0 = mems_0_0_io_rdata;
  assign FF_io_in = _T_159[3:0];
  assign FF_clock = clock;
  assign FF_reset = reset;
endmodule
module FIFOWidthConvert(
  input         clock,
  input         reset,
  input  [31:0] io_enq_0,
  input  [31:0] io_enq_1,
  input  [31:0] io_enq_2,
  input  [31:0] io_enq_3,
  input  [31:0] io_enq_4,
  input  [31:0] io_enq_5,
  input  [31:0] io_enq_6,
  input  [31:0] io_enq_7,
  input  [31:0] io_enq_8,
  input  [31:0] io_enq_9,
  input  [31:0] io_enq_10,
  input  [31:0] io_enq_11,
  input  [31:0] io_enq_12,
  input  [31:0] io_enq_13,
  input  [31:0] io_enq_14,
  input  [31:0] io_enq_15,
  input         io_enqVld,
  output [31:0] io_deq_0,
  output [31:0] io_deq_1,
  output [31:0] io_deq_2,
  output [31:0] io_deq_3,
  output [31:0] io_deq_4,
  output [31:0] io_deq_5,
  output [31:0] io_deq_6,
  output [31:0] io_deq_7,
  output [31:0] io_deq_8,
  output [31:0] io_deq_9,
  output [31:0] io_deq_10,
  output [31:0] io_deq_11,
  output [31:0] io_deq_12,
  output [31:0] io_deq_13,
  output [31:0] io_deq_14,
  output [31:0] io_deq_15,
  input         io_deqVld,
  output        io_full,
  output        io_empty,
  output        io_almostEmpty,
  output        io_almostFull
);
  wire  FIFOCore_clock;
  wire  FIFOCore_reset;
  wire [31:0] FIFOCore_io_enq_0;
  wire [31:0] FIFOCore_io_enq_1;
  wire [31:0] FIFOCore_io_enq_2;
  wire [31:0] FIFOCore_io_enq_3;
  wire [31:0] FIFOCore_io_enq_4;
  wire [31:0] FIFOCore_io_enq_5;
  wire [31:0] FIFOCore_io_enq_6;
  wire [31:0] FIFOCore_io_enq_7;
  wire [31:0] FIFOCore_io_enq_8;
  wire [31:0] FIFOCore_io_enq_9;
  wire [31:0] FIFOCore_io_enq_10;
  wire [31:0] FIFOCore_io_enq_11;
  wire [31:0] FIFOCore_io_enq_12;
  wire [31:0] FIFOCore_io_enq_13;
  wire [31:0] FIFOCore_io_enq_14;
  wire [31:0] FIFOCore_io_enq_15;
  wire  FIFOCore_io_enqVld;
  wire [31:0] FIFOCore_io_deq_0;
  wire [31:0] FIFOCore_io_deq_1;
  wire [31:0] FIFOCore_io_deq_2;
  wire [31:0] FIFOCore_io_deq_3;
  wire [31:0] FIFOCore_io_deq_4;
  wire [31:0] FIFOCore_io_deq_5;
  wire [31:0] FIFOCore_io_deq_6;
  wire [31:0] FIFOCore_io_deq_7;
  wire [31:0] FIFOCore_io_deq_8;
  wire [31:0] FIFOCore_io_deq_9;
  wire [31:0] FIFOCore_io_deq_10;
  wire [31:0] FIFOCore_io_deq_11;
  wire [31:0] FIFOCore_io_deq_12;
  wire [31:0] FIFOCore_io_deq_13;
  wire [31:0] FIFOCore_io_deq_14;
  wire [31:0] FIFOCore_io_deq_15;
  wire  FIFOCore_io_deqVld;
  wire  FIFOCore_io_full;
  wire  FIFOCore_io_empty;
  wire  FIFOCore_io_almostFull;
  wire  FIFOCore_io_almostEmpty;
  FIFOCore_2 FIFOCore (
    .clock(FIFOCore_clock),
    .reset(FIFOCore_reset),
    .io_enq_0(FIFOCore_io_enq_0),
    .io_enq_1(FIFOCore_io_enq_1),
    .io_enq_2(FIFOCore_io_enq_2),
    .io_enq_3(FIFOCore_io_enq_3),
    .io_enq_4(FIFOCore_io_enq_4),
    .io_enq_5(FIFOCore_io_enq_5),
    .io_enq_6(FIFOCore_io_enq_6),
    .io_enq_7(FIFOCore_io_enq_7),
    .io_enq_8(FIFOCore_io_enq_8),
    .io_enq_9(FIFOCore_io_enq_9),
    .io_enq_10(FIFOCore_io_enq_10),
    .io_enq_11(FIFOCore_io_enq_11),
    .io_enq_12(FIFOCore_io_enq_12),
    .io_enq_13(FIFOCore_io_enq_13),
    .io_enq_14(FIFOCore_io_enq_14),
    .io_enq_15(FIFOCore_io_enq_15),
    .io_enqVld(FIFOCore_io_enqVld),
    .io_deq_0(FIFOCore_io_deq_0),
    .io_deq_1(FIFOCore_io_deq_1),
    .io_deq_2(FIFOCore_io_deq_2),
    .io_deq_3(FIFOCore_io_deq_3),
    .io_deq_4(FIFOCore_io_deq_4),
    .io_deq_5(FIFOCore_io_deq_5),
    .io_deq_6(FIFOCore_io_deq_6),
    .io_deq_7(FIFOCore_io_deq_7),
    .io_deq_8(FIFOCore_io_deq_8),
    .io_deq_9(FIFOCore_io_deq_9),
    .io_deq_10(FIFOCore_io_deq_10),
    .io_deq_11(FIFOCore_io_deq_11),
    .io_deq_12(FIFOCore_io_deq_12),
    .io_deq_13(FIFOCore_io_deq_13),
    .io_deq_14(FIFOCore_io_deq_14),
    .io_deq_15(FIFOCore_io_deq_15),
    .io_deqVld(FIFOCore_io_deqVld),
    .io_full(FIFOCore_io_full),
    .io_empty(FIFOCore_io_empty),
    .io_almostFull(FIFOCore_io_almostFull),
    .io_almostEmpty(FIFOCore_io_almostEmpty)
  );
  assign io_deq_0 = FIFOCore_io_deq_0;
  assign io_deq_1 = FIFOCore_io_deq_1;
  assign io_deq_2 = FIFOCore_io_deq_2;
  assign io_deq_3 = FIFOCore_io_deq_3;
  assign io_deq_4 = FIFOCore_io_deq_4;
  assign io_deq_5 = FIFOCore_io_deq_5;
  assign io_deq_6 = FIFOCore_io_deq_6;
  assign io_deq_7 = FIFOCore_io_deq_7;
  assign io_deq_8 = FIFOCore_io_deq_8;
  assign io_deq_9 = FIFOCore_io_deq_9;
  assign io_deq_10 = FIFOCore_io_deq_10;
  assign io_deq_11 = FIFOCore_io_deq_11;
  assign io_deq_12 = FIFOCore_io_deq_12;
  assign io_deq_13 = FIFOCore_io_deq_13;
  assign io_deq_14 = FIFOCore_io_deq_14;
  assign io_deq_15 = FIFOCore_io_deq_15;
  assign io_full = FIFOCore_io_full;
  assign io_empty = FIFOCore_io_empty;
  assign io_almostEmpty = FIFOCore_io_almostEmpty;
  assign io_almostFull = FIFOCore_io_almostFull;
  assign FIFOCore_io_enq_0 = io_enq_0;
  assign FIFOCore_io_enq_1 = io_enq_1;
  assign FIFOCore_io_enq_2 = io_enq_2;
  assign FIFOCore_io_enq_3 = io_enq_3;
  assign FIFOCore_io_enq_4 = io_enq_4;
  assign FIFOCore_io_enq_5 = io_enq_5;
  assign FIFOCore_io_enq_6 = io_enq_6;
  assign FIFOCore_io_enq_7 = io_enq_7;
  assign FIFOCore_io_enq_8 = io_enq_8;
  assign FIFOCore_io_enq_9 = io_enq_9;
  assign FIFOCore_io_enq_10 = io_enq_10;
  assign FIFOCore_io_enq_11 = io_enq_11;
  assign FIFOCore_io_enq_12 = io_enq_12;
  assign FIFOCore_io_enq_13 = io_enq_13;
  assign FIFOCore_io_enq_14 = io_enq_14;
  assign FIFOCore_io_enq_15 = io_enq_15;
  assign FIFOCore_io_enqVld = io_enqVld;
  assign FIFOCore_io_deqVld = io_deqVld;
  assign FIFOCore_clock = clock;
  assign FIFOCore_reset = reset;
endmodule
module RetimeWrapper_51(
  input          clock,
  input          reset,
  input  [511:0] io_in,
  output [511:0] io_out
);
  wire [511:0] sr_out;
  wire [511:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(512), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FFType_47(
  input          clock,
  input          reset,
  input  [511:0] io_in,
  input  [511:0] io_init,
  output [511:0] io_out,
  input          io_enable
);
  wire [511:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [511:0] RetimeWrapper_io_in;
  wire [511:0] RetimeWrapper_io_out;
  wire [511:0] _T_10;
  wire [511:0] _GEN_0;
  wire [511:0] _GEN_1;
  RetimeWrapper_51 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? io_init : _T_10;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_10;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_10 = RetimeWrapper_io_out;
endmodule
module FF_49(
  input          clock,
  input          reset,
  input  [511:0] io_in,
  input  [511:0] io_init,
  output [511:0] io_out,
  input          io_enable
);
  wire  ff_clock;
  wire  ff_reset;
  wire [511:0] ff_io_in;
  wire [511:0] ff_io_init;
  wire [511:0] ff_io_out;
  wire  ff_io_enable;
  FFType_47 ff (
    .clock(ff_clock),
    .reset(ff_reset),
    .io_in(ff_io_in),
    .io_init(ff_io_init),
    .io_out(ff_io_out),
    .io_enable(ff_io_enable)
  );
  assign io_out = ff_io_out;
  assign ff_io_in = io_in;
  assign ff_io_init = io_init;
  assign ff_io_enable = io_enable;
  assign ff_clock = clock;
  assign ff_reset = reset;
endmodule
module FIFOCounter(
  input   clock,
  input   reset,
  input   io_enqVld,
  output  io_full
);
  wire  sizeUDC_clock;
  wire  sizeUDC_reset;
  wire [9:0] sizeUDC_io_strideInc;
  wire [9:0] sizeUDC_io_strideDec;
  wire  sizeUDC_io_inc;
  wire  sizeUDC_io_dec;
  wire [9:0] sizeUDC_io_out;
  wire [9:0] sizeUDC_io_nextInc;
  wire [9:0] sizeUDC_io_nextDec;
  wire [10:0] _T_21;
  wire [10:0] _T_22;
  wire [9:0] remainingSlots;
  wire  full;
  wire  _T_34;
  wire  writeEn;
  UpDownCtr sizeUDC (
    .clock(sizeUDC_clock),
    .reset(sizeUDC_reset),
    .io_strideInc(sizeUDC_io_strideInc),
    .io_strideDec(sizeUDC_io_strideDec),
    .io_inc(sizeUDC_io_inc),
    .io_dec(sizeUDC_io_dec),
    .io_out(sizeUDC_io_out),
    .io_nextInc(sizeUDC_io_nextInc),
    .io_nextDec(sizeUDC_io_nextDec)
  );
  assign _T_21 = 10'h200 - sizeUDC_io_out;
  assign _T_22 = $unsigned(_T_21);
  assign remainingSlots = _T_22[9:0];
  assign full = remainingSlots < 10'h1;
  assign _T_34 = ~ full;
  assign writeEn = io_enqVld & _T_34;
  assign io_full = full;
  assign sizeUDC_io_strideInc = 10'h1;
  assign sizeUDC_io_strideDec = 10'h1;
  assign sizeUDC_io_inc = writeEn;
  assign sizeUDC_io_dec = 1'h0;
  assign sizeUDC_clock = clock;
  assign sizeUDC_reset = reset;
endmodule
module MAGCore(
  input         clock,
  input         reset,
  input         io_enable,
  input         io_dram_cmd_ready,
  output        io_dram_cmd_valid,
  output [63:0] io_dram_cmd_bits_addr,
  output [31:0] io_dram_cmd_bits_size,
  output        io_dram_cmd_bits_isWr,
  output [25:0] io_dram_cmd_bits_tag_uid,
  output [5:0]  io_dram_cmd_bits_tag_streamId,
  input         io_dram_wdata_ready,
  output        io_dram_wdata_valid,
  output [31:0] io_dram_wdata_bits_wdata_0,
  output [31:0] io_dram_wdata_bits_wdata_1,
  output [31:0] io_dram_wdata_bits_wdata_2,
  output [31:0] io_dram_wdata_bits_wdata_3,
  output [31:0] io_dram_wdata_bits_wdata_4,
  output [31:0] io_dram_wdata_bits_wdata_5,
  output [31:0] io_dram_wdata_bits_wdata_6,
  output [31:0] io_dram_wdata_bits_wdata_7,
  output [31:0] io_dram_wdata_bits_wdata_8,
  output [31:0] io_dram_wdata_bits_wdata_9,
  output [31:0] io_dram_wdata_bits_wdata_10,
  output [31:0] io_dram_wdata_bits_wdata_11,
  output [31:0] io_dram_wdata_bits_wdata_12,
  output [31:0] io_dram_wdata_bits_wdata_13,
  output [31:0] io_dram_wdata_bits_wdata_14,
  output [31:0] io_dram_wdata_bits_wdata_15,
  output        io_dram_wdata_bits_wlast,
  output        io_dram_rresp_ready,
  input         io_dram_rresp_valid,
  input  [31:0] io_dram_rresp_bits_rdata_0,
  input  [31:0] io_dram_rresp_bits_rdata_1,
  input  [31:0] io_dram_rresp_bits_rdata_2,
  input  [31:0] io_dram_rresp_bits_rdata_3,
  input  [31:0] io_dram_rresp_bits_rdata_4,
  input  [31:0] io_dram_rresp_bits_rdata_5,
  input  [31:0] io_dram_rresp_bits_rdata_6,
  input  [31:0] io_dram_rresp_bits_rdata_7,
  input  [31:0] io_dram_rresp_bits_rdata_8,
  input  [31:0] io_dram_rresp_bits_rdata_9,
  input  [31:0] io_dram_rresp_bits_rdata_10,
  input  [31:0] io_dram_rresp_bits_rdata_11,
  input  [31:0] io_dram_rresp_bits_rdata_12,
  input  [31:0] io_dram_rresp_bits_rdata_13,
  input  [31:0] io_dram_rresp_bits_rdata_14,
  input  [31:0] io_dram_rresp_bits_rdata_15,
  input  [5:0]  io_dram_rresp_bits_tag_streamId,
  output        io_dram_wresp_ready,
  input         io_dram_wresp_valid,
  input  [5:0]  io_dram_wresp_bits_tag_streamId,
  output [31:0] io_debugSignals_0,
  output [31:0] io_debugSignals_1,
  output [31:0] io_debugSignals_2,
  output [31:0] io_debugSignals_3,
  output [31:0] io_debugSignals_4,
  output [31:0] io_debugSignals_5,
  output [31:0] io_debugSignals_6,
  output [31:0] io_debugSignals_7,
  output [31:0] io_debugSignals_8,
  output [31:0] io_debugSignals_9,
  output [31:0] io_debugSignals_10,
  output [31:0] io_debugSignals_11,
  output [31:0] io_debugSignals_12,
  output [31:0] io_debugSignals_13,
  output [31:0] io_debugSignals_14,
  output [31:0] io_debugSignals_15,
  output [31:0] io_debugSignals_16,
  output [31:0] io_debugSignals_17,
  output [31:0] io_debugSignals_18,
  output [31:0] io_debugSignals_19,
  output [31:0] io_debugSignals_20,
  output [31:0] io_debugSignals_21,
  output [31:0] io_debugSignals_22,
  output [31:0] io_debugSignals_23,
  output [31:0] io_debugSignals_24,
  output [31:0] io_debugSignals_25,
  output [31:0] io_debugSignals_26,
  output [31:0] io_debugSignals_27,
  output [31:0] io_debugSignals_28,
  output [31:0] io_debugSignals_29,
  output [31:0] io_debugSignals_30,
  output [31:0] io_debugSignals_31,
  output [31:0] io_debugSignals_32,
  output [31:0] io_debugSignals_33,
  output [31:0] io_debugSignals_34,
  output [31:0] io_debugSignals_35,
  output [31:0] io_debugSignals_36,
  output [31:0] io_debugSignals_37,
  output [31:0] io_debugSignals_38,
  output [31:0] io_debugSignals_39,
  output [31:0] io_debugSignals_40,
  output [31:0] io_debugSignals_41,
  output [31:0] io_debugSignals_42,
  output [31:0] io_debugSignals_43,
  output [31:0] io_debugSignals_44,
  output [31:0] io_debugSignals_45,
  output [31:0] io_debugSignals_46,
  output [31:0] io_debugSignals_47,
  output [31:0] io_debugSignals_48,
  output [31:0] io_debugSignals_49,
  output [31:0] io_debugSignals_50,
  output [31:0] io_debugSignals_51,
  output [31:0] io_debugSignals_52,
  output [31:0] io_debugSignals_53,
  output [31:0] io_debugSignals_54,
  output [31:0] io_debugSignals_55,
  output [31:0] io_debugSignals_56,
  output [31:0] io_debugSignals_57,
  output [31:0] io_debugSignals_58,
  output [31:0] io_debugSignals_59,
  output [31:0] io_debugSignals_60,
  output [31:0] io_debugSignals_61,
  output [31:0] io_debugSignals_62,
  output [31:0] io_debugSignals_63,
  output [31:0] io_debugSignals_64,
  output [31:0] io_debugSignals_65,
  output [31:0] io_debugSignals_66,
  output [31:0] io_debugSignals_67,
  output [31:0] io_debugSignals_68,
  output [31:0] io_debugSignals_69,
  output [31:0] io_debugSignals_70,
  output [31:0] io_debugSignals_71,
  output [31:0] io_debugSignals_72,
  output [31:0] io_debugSignals_73,
  output [31:0] io_debugSignals_74,
  output [31:0] io_debugSignals_75,
  output [31:0] io_debugSignals_76,
  output [31:0] io_debugSignals_77,
  output [31:0] io_debugSignals_78,
  output [31:0] io_debugSignals_79,
  output [31:0] io_debugSignals_80,
  output [31:0] io_debugSignals_81,
  output [31:0] io_debugSignals_82,
  output [31:0] io_debugSignals_83,
  output [31:0] io_debugSignals_84,
  output [31:0] io_debugSignals_85,
  output [31:0] io_debugSignals_86,
  output [31:0] io_debugSignals_87,
  output [31:0] io_debugSignals_88,
  output [31:0] io_debugSignals_89,
  output [31:0] io_debugSignals_90,
  output [31:0] io_debugSignals_91,
  output [31:0] io_debugSignals_92,
  output [31:0] io_debugSignals_93,
  output [31:0] io_debugSignals_94,
  output [31:0] io_debugSignals_95,
  output [31:0] io_debugSignals_96,
  output [31:0] io_debugSignals_97,
  output [31:0] io_debugSignals_98,
  output [31:0] io_debugSignals_99,
  output [31:0] io_debugSignals_100,
  output [31:0] io_debugSignals_101,
  output [31:0] io_debugSignals_102,
  output [31:0] io_debugSignals_103,
  output [31:0] io_debugSignals_104,
  output [31:0] io_debugSignals_105,
  output [31:0] io_debugSignals_106,
  output [31:0] io_debugSignals_107,
  output [31:0] io_debugSignals_108,
  output [31:0] io_debugSignals_109,
  output [31:0] io_debugSignals_110,
  output [31:0] io_debugSignals_111,
  output [31:0] io_debugSignals_112,
  output [31:0] io_debugSignals_113
);
  wire  cmdArbiter_clock;
  wire  cmdArbiter_reset;
  wire [63:0] cmdArbiter_io_fifo_0_deq_0_addr;
  wire  cmdArbiter_io_fifo_0_deq_0_isWr;
  wire [15:0] cmdArbiter_io_fifo_0_deq_0_size;
  wire  cmdArbiter_io_fifo_0_deqVld;
  wire  cmdArbiter_io_fifo_0_empty;
  wire  cmdArbiter_io_fifo_0_almostEmpty;
  wire [63:0] cmdArbiter_io_fifo_1_deq_0_addr;
  wire  cmdArbiter_io_fifo_1_deq_0_isWr;
  wire [15:0] cmdArbiter_io_fifo_1_deq_0_size;
  wire  cmdArbiter_io_fifo_1_deqVld;
  wire  cmdArbiter_io_fifo_1_empty;
  wire [63:0] cmdArbiter_io_deq_0_addr;
  wire  cmdArbiter_io_deq_0_isWr;
  wire [15:0] cmdArbiter_io_deq_0_size;
  wire  cmdArbiter_io_deqVld;
  wire  cmdArbiter_io_empty;
  wire  cmdArbiter_io_tag;
  wire  cmdFifos_0_clock;
  wire  cmdFifos_0_reset;
  wire [63:0] cmdFifos_0_io_deq_0_addr;
  wire  cmdFifos_0_io_deq_0_isWr;
  wire [15:0] cmdFifos_0_io_deq_0_size;
  wire  cmdFifos_0_io_deqVld;
  wire  cmdFifos_0_io_empty;
  wire  cmdFifos_0_io_almostEmpty;
  wire  cmdFifos_1_clock;
  wire  cmdFifos_1_reset;
  wire [63:0] cmdFifos_1_io_deq_0_addr;
  wire  cmdFifos_1_io_deq_0_isWr;
  wire [15:0] cmdFifos_1_io_deq_0_size;
  wire  cmdFifos_1_io_deqVld;
  wire  cmdFifos_1_io_empty;
  wire  cmdFifos_1_io_almostEmpty;
  wire [63:0] cmdAddr_bits;
  wire  _T_918;
  wire  _T_919;
  wire  _T_920;
  wire  cmdRead;
  wire  cmdWrite;
  wire  burstCounter_clock;
  wire  burstCounter_reset;
  wire [31:0] burstCounter_io_max;
  wire [31:0] burstCounter_io_out;
  wire  burstCounter_io_enable;
  wire  burstCounter_io_done;
  wire  burstTagCounter_clock;
  wire  burstTagCounter_reset;
  wire [9:0] burstTagCounter_io_max;
  wire [9:0] burstTagCounter_io_out;
  wire [9:0] burstTagCounter_io_next;
  wire  burstTagCounter_io_enable;
  wire  burstTagCounter_io_done;
  wire  dramReadySeen;
  wire  rrespReadyMux_io_ins_0;
  wire  rrespReadyMux_io_out;
  wire  wdataMux_io_ins_0_valid;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_0;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_1;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_2;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_3;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_4;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_5;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_6;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_7;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_8;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_9;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_10;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_11;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_12;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_13;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_14;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_15;
  wire  wdataMux_io_ins_0_bits_wlast;
  wire  wdataMux_io_out_valid;
  wire [31:0] wdataMux_io_out_bits_wdata_0;
  wire [31:0] wdataMux_io_out_bits_wdata_1;
  wire [31:0] wdataMux_io_out_bits_wdata_2;
  wire [31:0] wdataMux_io_out_bits_wdata_3;
  wire [31:0] wdataMux_io_out_bits_wdata_4;
  wire [31:0] wdataMux_io_out_bits_wdata_5;
  wire [31:0] wdataMux_io_out_bits_wdata_6;
  wire [31:0] wdataMux_io_out_bits_wdata_7;
  wire [31:0] wdataMux_io_out_bits_wdata_8;
  wire [31:0] wdataMux_io_out_bits_wdata_9;
  wire [31:0] wdataMux_io_out_bits_wdata_10;
  wire [31:0] wdataMux_io_out_bits_wdata_11;
  wire [31:0] wdataMux_io_out_bits_wdata_12;
  wire [31:0] wdataMux_io_out_bits_wdata_13;
  wire [31:0] wdataMux_io_out_bits_wdata_14;
  wire [31:0] wdataMux_io_out_bits_wdata_15;
  wire  wdataMux_io_out_bits_wlast;
  wire [32:0] _T_935;
  wire [32:0] _T_936;
  wire [31:0] _T_937;
  wire  _T_938;
  wire  _T_939;
  wire  cmdDeqValidMux_io_ins_0;
  wire  cmdDeqValidMux_io_ins_1;
  wire  cmdDeqValidMux_io_sel;
  wire  cmdDeqValidMux_io_out;
  wire  dramCmdMux_io_ins_0_valid;
  wire [63:0] dramCmdMux_io_ins_0_bits_addr;
  wire [31:0] dramCmdMux_io_ins_0_bits_size;
  wire  dramCmdMux_io_ins_0_bits_isWr;
  wire [25:0] dramCmdMux_io_ins_0_bits_tag_uid;
  wire [5:0] dramCmdMux_io_ins_0_bits_tag_streamId;
  wire  dramCmdMux_io_ins_1_valid;
  wire [63:0] dramCmdMux_io_ins_1_bits_addr;
  wire [31:0] dramCmdMux_io_ins_1_bits_size;
  wire  dramCmdMux_io_ins_1_bits_isWr;
  wire [25:0] dramCmdMux_io_ins_1_bits_tag_uid;
  wire [5:0] dramCmdMux_io_ins_1_bits_tag_streamId;
  wire  dramCmdMux_io_sel;
  wire  dramCmdMux_io_out_valid;
  wire [63:0] dramCmdMux_io_out_bits_addr;
  wire [31:0] dramCmdMux_io_out_bits_size;
  wire  dramCmdMux_io_out_bits_isWr;
  wire [25:0] dramCmdMux_io_out_bits_tag_uid;
  wire [5:0] dramCmdMux_io_out_bits_tag_streamId;
  wire [57:0] _T_942;
  wire [63:0] _T_944;
  wire [5:0] _T_946_streamId;
  wire [15:0] _T_948_bits;
  wire [9:0] _T_949;
  wire [5:0] _T_950;
  wire  _T_952;
  wire [9:0] _GEN_0;
  wire [10:0] _T_953;
  wire [9:0] _T_954;
  wire  _T_955;
  wire  _T_956;
  wire  FF_clock;
  wire  FF_reset;
  wire [5:0] FF_io_in;
  wire [5:0] FF_io_init;
  wire [5:0] FF_io_out;
  wire  FF_io_enable;
  wire  FF_1_clock;
  wire  FF_1_reset;
  wire [63:0] FF_1_io_in;
  wire [63:0] FF_1_io_init;
  wire [63:0] FF_1_io_out;
  wire  FF_1_io_enable;
  wire  FF_2_clock;
  wire  FF_2_reset;
  wire [31:0] FF_2_io_in;
  wire [31:0] FF_2_io_init;
  wire [31:0] FF_2_io_out;
  wire  FF_2_io_enable;
  wire [5:0] _T_974_streamId;
  wire [15:0] _T_976_bits;
  wire [9:0] _T_977;
  wire [5:0] _T_978;
  wire  _T_980;
  wire [9:0] _GEN_1;
  wire [10:0] _T_981;
  wire [9:0] _T_982;
  wire  FF_3_clock;
  wire  FF_3_reset;
  wire  FF_3_io_in;
  wire  FF_3_io_init;
  wire  FF_3_io_out;
  wire  FF_3_io_enable;
  wire  FF_4_clock;
  wire  FF_4_reset;
  wire [63:0] FF_4_io_in;
  wire [63:0] FF_4_io_init;
  wire [63:0] FF_4_io_out;
  wire  FF_4_io_enable;
  wire  FF_5_clock;
  wire  FF_5_reset;
  wire [15:0] FF_5_io_in;
  wire [15:0] FF_5_io_out;
  wire  FF_5_io_enable;
  wire  wrespReadyMux_io_ins_0;
  wire  wrespReadyMux_io_out;
  wire  gatherLoadIssueMux_io_ins_0;
  wire  gatherLoadIssueMux_io_ins_1;
  wire  gatherLoadIssueMux_io_sel;
  wire  gatherLoadIssueMux_io_out;
  wire  gatherLoadIssue_clock;
  wire  gatherLoadIssue_reset;
  wire [31:0] gatherLoadIssue_io_max;
  wire [31:0] gatherLoadIssue_io_out;
  wire  gatherLoadIssue_io_enable;
  wire  gatherLoadIssue_io_done;
  wire  gatherLoadSkipMux_io_ins_0;
  wire  gatherLoadSkipMux_io_ins_1;
  wire  gatherLoadSkipMux_io_sel;
  wire  gatherLoadSkipMux_io_out;
  wire  gatherLoadSkip_clock;
  wire  gatherLoadSkip_reset;
  wire [31:0] gatherLoadSkip_io_max;
  wire [31:0] gatherLoadSkip_io_out;
  wire  gatherLoadSkip_io_enable;
  wire  gatherLoadSkip_io_done;
  wire  scatterLoadIssueMux_io_ins_0;
  wire  scatterLoadIssueMux_io_ins_1;
  wire  scatterLoadIssueMux_io_sel;
  wire  scatterLoadIssueMux_io_out;
  wire  scatterLoadIssue_clock;
  wire  scatterLoadIssue_reset;
  wire [31:0] scatterLoadIssue_io_max;
  wire [31:0] scatterLoadIssue_io_out;
  wire  scatterLoadIssue_io_enable;
  wire  scatterLoadIssue_io_done;
  wire  scatterLoadSkipMux_io_ins_0;
  wire  scatterLoadSkipMux_io_ins_1;
  wire  scatterLoadSkipMux_io_sel;
  wire  scatterLoadSkipMux_io_out;
  wire  scatterLoadSkip_clock;
  wire  scatterLoadSkip_reset;
  wire [31:0] scatterLoadSkip_io_max;
  wire [31:0] scatterLoadSkip_io_out;
  wire  scatterLoadSkip_io_enable;
  wire  scatterLoadSkip_io_done;
  wire  scatterStoreIssueMux_io_ins_0;
  wire  scatterStoreIssueMux_io_ins_1;
  wire  scatterStoreIssueMux_io_sel;
  wire  scatterStoreIssueMux_io_out;
  wire  scatterStoreIssue_clock;
  wire  scatterStoreIssue_reset;
  wire [31:0] scatterStoreIssue_io_max;
  wire [31:0] scatterStoreIssue_io_out;
  wire  scatterStoreIssue_io_enable;
  wire  scatterStoreIssue_io_done;
  wire  scatterStoreSkipMux_io_ins_0;
  wire  scatterStoreSkipMux_io_ins_1;
  wire  scatterStoreSkipMux_io_sel;
  wire  scatterStoreSkipMux_io_out;
  wire  scatterStoreSkip_clock;
  wire  scatterStoreSkip_reset;
  wire [31:0] scatterStoreSkip_io_max;
  wire [31:0] scatterStoreSkip_io_out;
  wire  scatterStoreSkip_io_enable;
  wire  scatterStoreSkip_io_done;
  wire  denseLoadBuffers_0_clock;
  wire  denseLoadBuffers_0_reset;
  wire [31:0] denseLoadBuffers_0_io_enq_0;
  wire [31:0] denseLoadBuffers_0_io_enq_1;
  wire [31:0] denseLoadBuffers_0_io_enq_2;
  wire [31:0] denseLoadBuffers_0_io_enq_3;
  wire [31:0] denseLoadBuffers_0_io_enq_4;
  wire [31:0] denseLoadBuffers_0_io_enq_5;
  wire [31:0] denseLoadBuffers_0_io_enq_6;
  wire [31:0] denseLoadBuffers_0_io_enq_7;
  wire [31:0] denseLoadBuffers_0_io_enq_8;
  wire [31:0] denseLoadBuffers_0_io_enq_9;
  wire [31:0] denseLoadBuffers_0_io_enq_10;
  wire [31:0] denseLoadBuffers_0_io_enq_11;
  wire [31:0] denseLoadBuffers_0_io_enq_12;
  wire [31:0] denseLoadBuffers_0_io_enq_13;
  wire [31:0] denseLoadBuffers_0_io_enq_14;
  wire [31:0] denseLoadBuffers_0_io_enq_15;
  wire  denseLoadBuffers_0_io_enqVld;
  wire [31:0] denseLoadBuffers_0_io_deq_0;
  wire [31:0] denseLoadBuffers_0_io_deq_1;
  wire [31:0] denseLoadBuffers_0_io_deq_2;
  wire [31:0] denseLoadBuffers_0_io_deq_3;
  wire [31:0] denseLoadBuffers_0_io_deq_4;
  wire [31:0] denseLoadBuffers_0_io_deq_5;
  wire [31:0] denseLoadBuffers_0_io_deq_6;
  wire [31:0] denseLoadBuffers_0_io_deq_7;
  wire [31:0] denseLoadBuffers_0_io_deq_8;
  wire [31:0] denseLoadBuffers_0_io_deq_9;
  wire [31:0] denseLoadBuffers_0_io_deq_10;
  wire [31:0] denseLoadBuffers_0_io_deq_11;
  wire [31:0] denseLoadBuffers_0_io_deq_12;
  wire [31:0] denseLoadBuffers_0_io_deq_13;
  wire [31:0] denseLoadBuffers_0_io_deq_14;
  wire [31:0] denseLoadBuffers_0_io_deq_15;
  wire  denseLoadBuffers_0_io_deqVld;
  wire  denseLoadBuffers_0_io_full;
  wire  denseLoadBuffers_0_io_empty;
  wire  denseLoadBuffers_0_io_almostEmpty;
  wire  denseLoadBuffers_0_io_almostFull;
  wire  _T_1035;
  wire  _T_1036;
  wire  _T_1037;
  wire  Counter_clock;
  wire  Counter_reset;
  wire [31:0] Counter_io_max;
  wire [31:0] Counter_io_out;
  wire  Counter_io_enable;
  wire  Counter_io_done;
  wire  _T_1044;
  wire  Counter_1_clock;
  wire  Counter_1_reset;
  wire [31:0] Counter_1_io_max;
  wire [31:0] Counter_1_io_out;
  wire  Counter_1_io_enable;
  wire  Counter_1_io_done;
  wire  SRFF_sp_clock;
  wire  SRFF_sp_reset;
  wire  SRFF_sp_io_input_set;
  wire  SRFF_sp_io_input_reset;
  wire  SRFF_sp_io_input_asyn_reset;
  wire  SRFF_sp_io_output_data;
  wire  SRFF_sp_1_clock;
  wire  SRFF_sp_1_reset;
  wire  SRFF_sp_1_io_input_set;
  wire  SRFF_sp_1_io_input_reset;
  wire  SRFF_sp_1_io_input_asyn_reset;
  wire  SRFF_sp_1_io_output_data;
  wire  _T_1054;
  wire  _T_1055;
  reg  _T_1058;
  reg [31:0] _RAND_0;
  wire  _T_1064;
  wire  _T_1065;
  wire [63:0] _T_1066;
  wire [95:0] _T_1067;
  wire [127:0] _T_1068;
  wire [159:0] _T_1069;
  wire [191:0] _T_1070;
  wire [223:0] _T_1071;
  wire [255:0] _T_1072;
  wire [287:0] _T_1073;
  wire [319:0] _T_1074;
  wire [351:0] _T_1075;
  wire [383:0] _T_1076;
  wire [415:0] _T_1077;
  wire [447:0] _T_1078;
  wire [479:0] _T_1079;
  wire [511:0] _T_1080;
  wire  FF_6_clock;
  wire  FF_6_reset;
  wire [511:0] FF_6_io_in;
  wire [511:0] FF_6_io_init;
  wire [511:0] FF_6_io_out;
  wire  FF_6_io_enable;
  wire  _T_1084;
  wire  _T_1085;
  reg  _T_1088;
  reg [31:0] _RAND_1;
  wire  _T_1094;
  wire  _T_1095;
  wire [63:0] _T_1096;
  wire [95:0] _T_1097;
  wire [127:0] _T_1098;
  wire [159:0] _T_1099;
  wire [191:0] _T_1100;
  wire [223:0] _T_1101;
  wire [255:0] _T_1102;
  wire [287:0] _T_1103;
  wire [319:0] _T_1104;
  wire [351:0] _T_1105;
  wire [383:0] _T_1106;
  wire [415:0] _T_1107;
  wire [447:0] _T_1108;
  wire [479:0] _T_1109;
  wire [511:0] _T_1110;
  wire  FF_7_clock;
  wire  FF_7_reset;
  wire [511:0] FF_7_io_in;
  wire [511:0] FF_7_io_init;
  wire [511:0] FF_7_io_out;
  wire  FF_7_io_enable;
  wire  denseStoreBuffers_0_clock;
  wire  denseStoreBuffers_0_reset;
  wire [31:0] denseStoreBuffers_0_io_enq_0;
  wire [31:0] denseStoreBuffers_0_io_enq_1;
  wire [31:0] denseStoreBuffers_0_io_enq_2;
  wire [31:0] denseStoreBuffers_0_io_enq_3;
  wire [31:0] denseStoreBuffers_0_io_enq_4;
  wire [31:0] denseStoreBuffers_0_io_enq_5;
  wire [31:0] denseStoreBuffers_0_io_enq_6;
  wire [31:0] denseStoreBuffers_0_io_enq_7;
  wire [31:0] denseStoreBuffers_0_io_enq_8;
  wire [31:0] denseStoreBuffers_0_io_enq_9;
  wire [31:0] denseStoreBuffers_0_io_enq_10;
  wire [31:0] denseStoreBuffers_0_io_enq_11;
  wire [31:0] denseStoreBuffers_0_io_enq_12;
  wire [31:0] denseStoreBuffers_0_io_enq_13;
  wire [31:0] denseStoreBuffers_0_io_enq_14;
  wire [31:0] denseStoreBuffers_0_io_enq_15;
  wire  denseStoreBuffers_0_io_enqVld;
  wire [31:0] denseStoreBuffers_0_io_deq_0;
  wire [31:0] denseStoreBuffers_0_io_deq_1;
  wire [31:0] denseStoreBuffers_0_io_deq_2;
  wire [31:0] denseStoreBuffers_0_io_deq_3;
  wire [31:0] denseStoreBuffers_0_io_deq_4;
  wire [31:0] denseStoreBuffers_0_io_deq_5;
  wire [31:0] denseStoreBuffers_0_io_deq_6;
  wire [31:0] denseStoreBuffers_0_io_deq_7;
  wire [31:0] denseStoreBuffers_0_io_deq_8;
  wire [31:0] denseStoreBuffers_0_io_deq_9;
  wire [31:0] denseStoreBuffers_0_io_deq_10;
  wire [31:0] denseStoreBuffers_0_io_deq_11;
  wire [31:0] denseStoreBuffers_0_io_deq_12;
  wire [31:0] denseStoreBuffers_0_io_deq_13;
  wire [31:0] denseStoreBuffers_0_io_deq_14;
  wire [31:0] denseStoreBuffers_0_io_deq_15;
  wire  denseStoreBuffers_0_io_deqVld;
  wire  denseStoreBuffers_0_io_full;
  wire  denseStoreBuffers_0_io_empty;
  wire  denseStoreBuffers_0_io_almostEmpty;
  wire  denseStoreBuffers_0_io_almostFull;
  wire  _T_1114;
  wire  _T_1115;
  wire  _T_1116;
  wire  _T_1117;
  wire  _T_1118;
  wire  _T_1119;
  wire  _T_1121;
  wire  _T_1122;
  wire  FIFOCounter_clock;
  wire  FIFOCounter_reset;
  wire  FIFOCounter_io_enqVld;
  wire  FIFOCounter_io_full;
  wire  _T_1127;
  wire  _T_1128;
  wire  _T_1129;
  wire  Counter_2_clock;
  wire  Counter_2_reset;
  wire [31:0] Counter_2_io_max;
  wire [31:0] Counter_2_io_out;
  wire  Counter_2_io_enable;
  wire  Counter_2_io_done;
  wire [31:0] _T_1137;
  wire  _T_1140;
  wire  _T_1141;
  wire  _T_1142;
  wire  dramReadyFF_clock;
  wire  dramReadyFF_reset;
  wire  dramReadyFF_io_in;
  wire  dramReadyFF_io_init;
  wire  dramReadyFF_io_out;
  wire  dramReadyFF_io_enable;
  wire  _T_1150;
  wire  _T_1151;
  wire  _T_1153;
  wire  _T_1154;
  wire  cycleCount_clock;
  wire  cycleCount_reset;
  wire [31:0] cycleCount_io_max;
  wire [31:0] cycleCount_io_out;
  wire  cycleCount_io_enable;
  wire  cycleCount_io_done;
  wire  _T_1160;
  wire  rdataEnqCount_clock;
  wire  rdataEnqCount_reset;
  wire [31:0] rdataEnqCount_io_max;
  wire [31:0] rdataEnqCount_io_out;
  wire  rdataEnqCount_io_enable;
  wire  rdataEnqCount_io_done;
  wire  _T_1166;
  wire  _T_1167;
  wire  wdataCount_clock;
  wire  wdataCount_reset;
  wire [31:0] wdataCount_io_max;
  wire [31:0] wdataCount_io_out;
  wire  wdataCount_io_enable;
  wire  wdataCount_io_done;
  wire  _T_1173;
  wire  _T_1175;
  wire  _T_1176;
  wire  FF_8_clock;
  wire  FF_8_reset;
  wire [31:0] FF_8_io_in;
  wire [31:0] FF_8_io_init;
  wire [31:0] FF_8_io_out;
  wire  FF_8_io_enable;
  wire  FF_9_clock;
  wire  FF_9_reset;
  wire [31:0] FF_9_io_in;
  wire [31:0] FF_9_io_init;
  wire [31:0] FF_9_io_out;
  wire  FF_9_io_enable;
  wire  FF_10_clock;
  wire  FF_10_reset;
  wire [31:0] FF_10_io_in;
  wire [31:0] FF_10_io_init;
  wire [31:0] FF_10_io_out;
  wire  FF_10_io_enable;
  wire  FF_11_clock;
  wire  FF_11_reset;
  wire [31:0] FF_11_io_in;
  wire [31:0] FF_11_io_init;
  wire [31:0] FF_11_io_out;
  wire  FF_11_io_enable;
  wire  FF_12_clock;
  wire  FF_12_reset;
  wire [31:0] FF_12_io_in;
  wire [31:0] FF_12_io_init;
  wire [31:0] FF_12_io_out;
  wire  FF_12_io_enable;
  wire  FF_13_clock;
  wire  FF_13_reset;
  wire [31:0] FF_13_io_in;
  wire [31:0] FF_13_io_init;
  wire [31:0] FF_13_io_out;
  wire  FF_13_io_enable;
  wire  FF_14_clock;
  wire  FF_14_reset;
  wire [31:0] FF_14_io_in;
  wire [31:0] FF_14_io_init;
  wire [31:0] FF_14_io_out;
  wire  FF_14_io_enable;
  wire  FF_15_clock;
  wire  FF_15_reset;
  wire [31:0] FF_15_io_in;
  wire [31:0] FF_15_io_init;
  wire [31:0] FF_15_io_out;
  wire  FF_15_io_enable;
  wire  FF_16_clock;
  wire  FF_16_reset;
  wire [31:0] FF_16_io_in;
  wire [31:0] FF_16_io_init;
  wire [31:0] FF_16_io_out;
  wire  FF_16_io_enable;
  wire  FF_17_clock;
  wire  FF_17_reset;
  wire [31:0] FF_17_io_in;
  wire [31:0] FF_17_io_init;
  wire [31:0] FF_17_io_out;
  wire  FF_17_io_enable;
  wire  FF_18_clock;
  wire  FF_18_reset;
  wire [31:0] FF_18_io_in;
  wire [31:0] FF_18_io_init;
  wire [31:0] FF_18_io_out;
  wire  FF_18_io_enable;
  wire  FF_19_clock;
  wire  FF_19_reset;
  wire [31:0] FF_19_io_in;
  wire [31:0] FF_19_io_init;
  wire [31:0] FF_19_io_out;
  wire  FF_19_io_enable;
  wire  FF_20_clock;
  wire  FF_20_reset;
  wire [31:0] FF_20_io_in;
  wire [31:0] FF_20_io_init;
  wire [31:0] FF_20_io_out;
  wire  FF_20_io_enable;
  wire  FF_21_clock;
  wire  FF_21_reset;
  wire [31:0] FF_21_io_in;
  wire [31:0] FF_21_io_init;
  wire [31:0] FF_21_io_out;
  wire  FF_21_io_enable;
  wire  FF_22_clock;
  wire  FF_22_reset;
  wire [31:0] FF_22_io_in;
  wire [31:0] FF_22_io_init;
  wire [31:0] FF_22_io_out;
  wire  FF_22_io_enable;
  wire  FF_23_clock;
  wire  FF_23_reset;
  wire [31:0] FF_23_io_in;
  wire [31:0] FF_23_io_init;
  wire [31:0] FF_23_io_out;
  wire  FF_23_io_enable;
  wire  _T_1287;
  wire  _T_1288;
  wire  FF_24_clock;
  wire  FF_24_reset;
  wire [31:0] FF_24_io_in;
  wire [31:0] FF_24_io_init;
  wire [31:0] FF_24_io_out;
  wire  FF_24_io_enable;
  wire  FF_25_clock;
  wire  FF_25_reset;
  wire [31:0] FF_25_io_in;
  wire [31:0] FF_25_io_init;
  wire [31:0] FF_25_io_out;
  wire  FF_25_io_enable;
  wire  FF_26_clock;
  wire  FF_26_reset;
  wire [31:0] FF_26_io_in;
  wire [31:0] FF_26_io_init;
  wire [31:0] FF_26_io_out;
  wire  FF_26_io_enable;
  wire  FF_27_clock;
  wire  FF_27_reset;
  wire [31:0] FF_27_io_in;
  wire [31:0] FF_27_io_init;
  wire [31:0] FF_27_io_out;
  wire  FF_27_io_enable;
  wire  FF_28_clock;
  wire  FF_28_reset;
  wire [31:0] FF_28_io_in;
  wire [31:0] FF_28_io_init;
  wire [31:0] FF_28_io_out;
  wire  FF_28_io_enable;
  wire  FF_29_clock;
  wire  FF_29_reset;
  wire [31:0] FF_29_io_in;
  wire [31:0] FF_29_io_init;
  wire [31:0] FF_29_io_out;
  wire  FF_29_io_enable;
  wire  FF_30_clock;
  wire  FF_30_reset;
  wire [31:0] FF_30_io_in;
  wire [31:0] FF_30_io_init;
  wire [31:0] FF_30_io_out;
  wire  FF_30_io_enable;
  wire  FF_31_clock;
  wire  FF_31_reset;
  wire [31:0] FF_31_io_in;
  wire [31:0] FF_31_io_init;
  wire [31:0] FF_31_io_out;
  wire  FF_31_io_enable;
  wire  FF_32_clock;
  wire  FF_32_reset;
  wire [31:0] FF_32_io_in;
  wire [31:0] FF_32_io_init;
  wire [31:0] FF_32_io_out;
  wire  FF_32_io_enable;
  wire  FF_33_clock;
  wire  FF_33_reset;
  wire [31:0] FF_33_io_in;
  wire [31:0] FF_33_io_init;
  wire [31:0] FF_33_io_out;
  wire  FF_33_io_enable;
  wire  FF_34_clock;
  wire  FF_34_reset;
  wire [31:0] FF_34_io_in;
  wire [31:0] FF_34_io_init;
  wire [31:0] FF_34_io_out;
  wire  FF_34_io_enable;
  wire  FF_35_clock;
  wire  FF_35_reset;
  wire [31:0] FF_35_io_in;
  wire [31:0] FF_35_io_init;
  wire [31:0] FF_35_io_out;
  wire  FF_35_io_enable;
  wire  FF_36_clock;
  wire  FF_36_reset;
  wire [31:0] FF_36_io_in;
  wire [31:0] FF_36_io_init;
  wire [31:0] FF_36_io_out;
  wire  FF_36_io_enable;
  wire  FF_37_clock;
  wire  FF_37_reset;
  wire [31:0] FF_37_io_in;
  wire [31:0] FF_37_io_init;
  wire [31:0] FF_37_io_out;
  wire  FF_37_io_enable;
  wire  FF_38_clock;
  wire  FF_38_reset;
  wire [31:0] FF_38_io_in;
  wire [31:0] FF_38_io_init;
  wire [31:0] FF_38_io_out;
  wire  FF_38_io_enable;
  wire  FF_39_clock;
  wire  FF_39_reset;
  wire [31:0] FF_39_io_in;
  wire [31:0] FF_39_io_init;
  wire [31:0] FF_39_io_out;
  wire  FF_39_io_enable;
  wire  _T_1397;
  wire  _T_1399;
  wire  _T_1400;
  wire  FF_40_clock;
  wire  FF_40_reset;
  wire [31:0] FF_40_io_in;
  wire [31:0] FF_40_io_init;
  wire [31:0] FF_40_io_out;
  wire  FF_40_io_enable;
  wire  FF_41_clock;
  wire  FF_41_reset;
  wire [31:0] FF_41_io_in;
  wire [31:0] FF_41_io_init;
  wire [31:0] FF_41_io_out;
  wire  FF_41_io_enable;
  wire  FF_42_clock;
  wire  FF_42_reset;
  wire [31:0] FF_42_io_in;
  wire [31:0] FF_42_io_init;
  wire [31:0] FF_42_io_out;
  wire  FF_42_io_enable;
  wire  FF_43_clock;
  wire  FF_43_reset;
  wire [31:0] FF_43_io_in;
  wire [31:0] FF_43_io_init;
  wire [31:0] FF_43_io_out;
  wire  FF_43_io_enable;
  wire  FF_44_clock;
  wire  FF_44_reset;
  wire [31:0] FF_44_io_in;
  wire [31:0] FF_44_io_init;
  wire [31:0] FF_44_io_out;
  wire  FF_44_io_enable;
  wire  FF_45_clock;
  wire  FF_45_reset;
  wire [31:0] FF_45_io_in;
  wire [31:0] FF_45_io_init;
  wire [31:0] FF_45_io_out;
  wire  FF_45_io_enable;
  wire  FF_46_clock;
  wire  FF_46_reset;
  wire [31:0] FF_46_io_in;
  wire [31:0] FF_46_io_init;
  wire [31:0] FF_46_io_out;
  wire  FF_46_io_enable;
  wire  FF_47_clock;
  wire  FF_47_reset;
  wire [31:0] FF_47_io_in;
  wire [31:0] FF_47_io_init;
  wire [31:0] FF_47_io_out;
  wire  FF_47_io_enable;
  wire  FF_48_clock;
  wire  FF_48_reset;
  wire [31:0] FF_48_io_in;
  wire [31:0] FF_48_io_init;
  wire [31:0] FF_48_io_out;
  wire  FF_48_io_enable;
  wire  FF_49_clock;
  wire  FF_49_reset;
  wire [31:0] FF_49_io_in;
  wire [31:0] FF_49_io_init;
  wire [31:0] FF_49_io_out;
  wire  FF_49_io_enable;
  wire  FF_50_clock;
  wire  FF_50_reset;
  wire [31:0] FF_50_io_in;
  wire [31:0] FF_50_io_init;
  wire [31:0] FF_50_io_out;
  wire  FF_50_io_enable;
  wire  FF_51_clock;
  wire  FF_51_reset;
  wire [31:0] FF_51_io_in;
  wire [31:0] FF_51_io_init;
  wire [31:0] FF_51_io_out;
  wire  FF_51_io_enable;
  wire  FF_52_clock;
  wire  FF_52_reset;
  wire [31:0] FF_52_io_in;
  wire [31:0] FF_52_io_init;
  wire [31:0] FF_52_io_out;
  wire  FF_52_io_enable;
  wire  FF_53_clock;
  wire  FF_53_reset;
  wire [31:0] FF_53_io_in;
  wire [31:0] FF_53_io_init;
  wire [31:0] FF_53_io_out;
  wire  FF_53_io_enable;
  wire  FF_54_clock;
  wire  FF_54_reset;
  wire [31:0] FF_54_io_in;
  wire [31:0] FF_54_io_init;
  wire [31:0] FF_54_io_out;
  wire  FF_54_io_enable;
  wire  FF_55_clock;
  wire  FF_55_reset;
  wire [31:0] FF_55_io_in;
  wire [31:0] FF_55_io_init;
  wire [31:0] FF_55_io_out;
  wire  FF_55_io_enable;
  wire [63:0] _T_1513;
  wire [95:0] _T_1514;
  wire [127:0] _T_1515;
  wire [159:0] _T_1516;
  wire [191:0] _T_1517;
  wire [223:0] _T_1518;
  wire [255:0] _T_1519;
  wire [287:0] _T_1520;
  wire [319:0] _T_1521;
  wire [351:0] _T_1522;
  wire [383:0] _T_1523;
  wire [415:0] _T_1524;
  wire [447:0] _T_1525;
  wire [479:0] _T_1526;
  wire [511:0] _T_1527;
  wire  FF_56_clock;
  wire  FF_56_reset;
  wire [511:0] FF_56_io_in;
  wire [511:0] FF_56_io_init;
  wire [511:0] FF_56_io_out;
  wire  FF_56_io_enable;
  wire  _T_1533;
  wire  _T_1534;
  wire  FF_57_clock;
  wire  FF_57_reset;
  wire [31:0] FF_57_io_in;
  wire [31:0] FF_57_io_init;
  wire [31:0] FF_57_io_out;
  wire  FF_57_io_enable;
  wire  FF_58_clock;
  wire  FF_58_reset;
  wire [31:0] FF_58_io_in;
  wire [31:0] FF_58_io_init;
  wire [31:0] FF_58_io_out;
  wire  FF_58_io_enable;
  wire  FF_59_clock;
  wire  FF_59_reset;
  wire [31:0] FF_59_io_in;
  wire [31:0] FF_59_io_init;
  wire [31:0] FF_59_io_out;
  wire  FF_59_io_enable;
  wire  FF_60_clock;
  wire  FF_60_reset;
  wire [31:0] FF_60_io_in;
  wire [31:0] FF_60_io_init;
  wire [31:0] FF_60_io_out;
  wire  FF_60_io_enable;
  wire  FF_61_clock;
  wire  FF_61_reset;
  wire [31:0] FF_61_io_in;
  wire [31:0] FF_61_io_init;
  wire [31:0] FF_61_io_out;
  wire  FF_61_io_enable;
  wire  FF_62_clock;
  wire  FF_62_reset;
  wire [31:0] FF_62_io_in;
  wire [31:0] FF_62_io_init;
  wire [31:0] FF_62_io_out;
  wire  FF_62_io_enable;
  wire  FF_63_clock;
  wire  FF_63_reset;
  wire [31:0] FF_63_io_in;
  wire [31:0] FF_63_io_init;
  wire [31:0] FF_63_io_out;
  wire  FF_63_io_enable;
  wire  FF_64_clock;
  wire  FF_64_reset;
  wire [31:0] FF_64_io_in;
  wire [31:0] FF_64_io_init;
  wire [31:0] FF_64_io_out;
  wire  FF_64_io_enable;
  wire  FF_65_clock;
  wire  FF_65_reset;
  wire [31:0] FF_65_io_in;
  wire [31:0] FF_65_io_init;
  wire [31:0] FF_65_io_out;
  wire  FF_65_io_enable;
  wire  FF_66_clock;
  wire  FF_66_reset;
  wire [31:0] FF_66_io_in;
  wire [31:0] FF_66_io_init;
  wire [31:0] FF_66_io_out;
  wire  FF_66_io_enable;
  wire  FF_67_clock;
  wire  FF_67_reset;
  wire [31:0] FF_67_io_in;
  wire [31:0] FF_67_io_init;
  wire [31:0] FF_67_io_out;
  wire  FF_67_io_enable;
  wire  FF_68_clock;
  wire  FF_68_reset;
  wire [31:0] FF_68_io_in;
  wire [31:0] FF_68_io_init;
  wire [31:0] FF_68_io_out;
  wire  FF_68_io_enable;
  wire  FF_69_clock;
  wire  FF_69_reset;
  wire [31:0] FF_69_io_in;
  wire [31:0] FF_69_io_init;
  wire [31:0] FF_69_io_out;
  wire  FF_69_io_enable;
  wire  FF_70_clock;
  wire  FF_70_reset;
  wire [31:0] FF_70_io_in;
  wire [31:0] FF_70_io_init;
  wire [31:0] FF_70_io_out;
  wire  FF_70_io_enable;
  wire  FF_71_clock;
  wire  FF_71_reset;
  wire [31:0] FF_71_io_in;
  wire [31:0] FF_71_io_init;
  wire [31:0] FF_71_io_out;
  wire  FF_71_io_enable;
  wire  FF_72_clock;
  wire  FF_72_reset;
  wire [31:0] FF_72_io_in;
  wire [31:0] FF_72_io_init;
  wire [31:0] FF_72_io_out;
  wire  FF_72_io_enable;
  wire  FF_73_clock;
  wire  FF_73_reset;
  wire [511:0] FF_73_io_in;
  wire [511:0] FF_73_io_init;
  wire [511:0] FF_73_io_out;
  wire  FF_73_io_enable;
  wire  _T_1665;
  wire  _T_1666;
  wire  Counter_3_clock;
  wire  Counter_3_reset;
  wire [31:0] Counter_3_io_max;
  wire [31:0] Counter_3_io_out;
  wire  Counter_3_io_enable;
  wire  Counter_3_io_done;
  wire  _T_1674;
  wire  _T_1675;
  wire  _T_1676;
  wire  Counter_4_clock;
  wire  Counter_4_reset;
  wire [31:0] Counter_4_io_max;
  wire [31:0] Counter_4_io_out;
  wire  Counter_4_io_enable;
  wire  Counter_4_io_done;
  wire  _T_1685;
  wire  Counter_5_clock;
  wire  Counter_5_reset;
  wire [31:0] Counter_5_io_max;
  wire [31:0] Counter_5_io_out;
  wire  Counter_5_io_enable;
  wire  Counter_5_io_done;
  wire  Counter_6_clock;
  wire  Counter_6_reset;
  wire [31:0] Counter_6_io_max;
  wire [31:0] Counter_6_io_out;
  wire  Counter_6_io_enable;
  wire  Counter_6_io_done;
  wire  Counter_7_clock;
  wire  Counter_7_reset;
  wire [31:0] Counter_7_io_max;
  wire [31:0] Counter_7_io_out;
  wire  Counter_7_io_enable;
  wire  Counter_7_io_done;
  wire  _T_1706;
  wire  _T_1707;
  wire  Counter_8_clock;
  wire  Counter_8_reset;
  wire [31:0] Counter_8_io_max;
  wire [31:0] Counter_8_io_out;
  wire  Counter_8_io_enable;
  wire  Counter_8_io_done;
  wire  _T_1715;
  wire  Counter_9_clock;
  wire  Counter_9_reset;
  wire [31:0] Counter_9_io_max;
  wire [31:0] Counter_9_io_out;
  wire  Counter_9_io_enable;
  wire  Counter_9_io_done;
  wire  Counter_10_clock;
  wire  Counter_10_reset;
  wire [31:0] Counter_10_io_max;
  wire [31:0] Counter_10_io_out;
  wire  Counter_10_io_enable;
  wire  Counter_10_io_done;
  wire  Counter_11_clock;
  wire  Counter_11_reset;
  wire [31:0] Counter_11_io_max;
  wire [31:0] Counter_11_io_out;
  wire  Counter_11_io_enable;
  wire  Counter_11_io_done;
  wire  _T_1737;
  wire  Counter_12_clock;
  wire  Counter_12_reset;
  wire [31:0] Counter_12_io_max;
  wire [31:0] Counter_12_io_out;
  wire  Counter_12_io_enable;
  wire  Counter_12_io_done;
  wire  Counter_13_clock;
  wire  Counter_13_reset;
  wire [31:0] Counter_13_io_max;
  wire [31:0] Counter_13_io_out;
  wire  Counter_13_io_enable;
  wire  Counter_13_io_done;
  wire  _T_1749;
  wire  _T_1750;
  wire  _T_1751;
  wire  Counter_14_clock;
  wire  Counter_14_reset;
  wire [31:0] Counter_14_io_max;
  wire [31:0] Counter_14_io_out;
  wire  Counter_14_io_enable;
  wire  Counter_14_io_done;
  wire  _T_1757;
  wire  _T_1758;
  wire  _T_1759;
  wire  Counter_15_clock;
  wire  Counter_15_reset;
  wire [31:0] Counter_15_io_max;
  wire [31:0] Counter_15_io_out;
  wire  Counter_15_io_enable;
  wire  Counter_15_io_done;
  wire  _T_1768;
  wire  Counter_16_clock;
  wire  Counter_16_reset;
  wire [31:0] Counter_16_io_max;
  wire [31:0] Counter_16_io_out;
  wire  Counter_16_io_enable;
  wire  Counter_16_io_done;
  wire  _T_1774;
  wire  Counter_17_clock;
  wire  Counter_17_reset;
  wire [31:0] Counter_17_io_max;
  wire [31:0] Counter_17_io_out;
  wire  Counter_17_io_enable;
  wire  Counter_17_io_done;
  wire  _T_1780;
  wire  _T_1781;
  wire  _T_1782;
  wire  Counter_18_clock;
  wire  Counter_18_reset;
  wire [31:0] Counter_18_io_max;
  wire [31:0] Counter_18_io_out;
  wire  Counter_18_io_enable;
  wire  Counter_18_io_done;
  wire  _T_1788;
  wire  _T_1789;
  wire  _T_1790;
  wire  Counter_19_clock;
  wire  Counter_19_reset;
  wire [31:0] Counter_19_io_max;
  wire [31:0] Counter_19_io_out;
  wire  Counter_19_io_enable;
  wire  Counter_19_io_done;
  wire  _T_1799;
  wire  Counter_20_clock;
  wire  Counter_20_reset;
  wire [31:0] Counter_20_io_max;
  wire [31:0] Counter_20_io_out;
  wire  Counter_20_io_enable;
  wire  Counter_20_io_done;
  wire  Counter_21_clock;
  wire  Counter_21_reset;
  wire [31:0] Counter_21_io_max;
  wire [31:0] Counter_21_io_out;
  wire  Counter_21_io_enable;
  wire  Counter_21_io_done;
  wire  Counter_22_clock;
  wire  Counter_22_reset;
  wire [31:0] Counter_22_io_max;
  wire [31:0] Counter_22_io_out;
  wire  Counter_22_io_enable;
  wire  Counter_22_io_done;
  wire  Counter_23_clock;
  wire  Counter_23_reset;
  wire [31:0] Counter_23_io_max;
  wire [31:0] Counter_23_io_out;
  wire  Counter_23_io_enable;
  wire  Counter_23_io_done;
  wire  Counter_24_clock;
  wire  Counter_24_reset;
  wire [31:0] Counter_24_io_max;
  wire [31:0] Counter_24_io_out;
  wire  Counter_24_io_enable;
  wire  Counter_24_io_done;
  wire  Counter_25_clock;
  wire  Counter_25_reset;
  wire [31:0] Counter_25_io_max;
  wire [31:0] Counter_25_io_out;
  wire  Counter_25_io_enable;
  wire  Counter_25_io_done;
  wire  Counter_26_clock;
  wire  Counter_26_reset;
  wire [31:0] Counter_26_io_max;
  wire [31:0] Counter_26_io_out;
  wire  Counter_26_io_enable;
  wire  Counter_26_io_done;
  wire  Counter_27_clock;
  wire  Counter_27_reset;
  wire [31:0] Counter_27_io_max;
  wire [31:0] Counter_27_io_out;
  wire  Counter_27_io_enable;
  wire  Counter_27_io_done;
  wire  _T_1843;
  wire  Counter_28_clock;
  wire  Counter_28_reset;
  wire [31:0] Counter_28_io_max;
  wire [31:0] Counter_28_io_out;
  wire  Counter_28_io_enable;
  wire  Counter_28_io_done;
  wire  FF_74_clock;
  wire  FF_74_reset;
  wire [5:0] FF_74_io_in;
  wire [5:0] FF_74_io_init;
  wire [5:0] FF_74_io_out;
  wire  FF_74_io_enable;
  wire  Counter_29_clock;
  wire  Counter_29_reset;
  wire [31:0] Counter_29_io_max;
  wire [31:0] Counter_29_io_out;
  wire  Counter_29_io_enable;
  wire  Counter_29_io_done;
  wire  Counter_30_clock;
  wire  Counter_30_reset;
  wire [31:0] Counter_30_io_max;
  wire [31:0] Counter_30_io_out;
  wire  Counter_30_io_enable;
  wire  Counter_30_io_done;
  wire  Counter_31_clock;
  wire  Counter_31_reset;
  wire [31:0] Counter_31_io_max;
  wire [31:0] Counter_31_io_out;
  wire  Counter_31_io_enable;
  wire  Counter_31_io_done;
  wire  Counter_32_clock;
  wire  Counter_32_reset;
  wire [31:0] Counter_32_io_max;
  wire [31:0] Counter_32_io_out;
  wire  Counter_32_io_enable;
  wire  Counter_32_io_done;
  wire  _T_1872;
  wire  Counter_33_clock;
  wire  Counter_33_reset;
  wire [31:0] Counter_33_io_max;
  wire [31:0] Counter_33_io_out;
  wire  Counter_33_io_enable;
  wire  Counter_33_io_done;
  wire  Counter_34_clock;
  wire  Counter_34_reset;
  wire [31:0] Counter_34_io_max;
  wire [31:0] Counter_34_io_out;
  wire  Counter_34_io_enable;
  wire  Counter_34_io_done;
  wire  _T_1885;
  wire  Counter_35_clock;
  wire  Counter_35_reset;
  wire [31:0] Counter_35_io_max;
  wire [31:0] Counter_35_io_out;
  wire  Counter_35_io_enable;
  wire  Counter_35_io_done;
  wire  _T_1892;
  wire  Counter_36_clock;
  wire  Counter_36_reset;
  wire [31:0] Counter_36_io_max;
  wire [31:0] Counter_36_io_out;
  wire  Counter_36_io_enable;
  wire  Counter_36_io_done;
  FIFOArbiter cmdArbiter (
    .clock(cmdArbiter_clock),
    .reset(cmdArbiter_reset),
    .io_fifo_0_deq_0_addr(cmdArbiter_io_fifo_0_deq_0_addr),
    .io_fifo_0_deq_0_isWr(cmdArbiter_io_fifo_0_deq_0_isWr),
    .io_fifo_0_deq_0_size(cmdArbiter_io_fifo_0_deq_0_size),
    .io_fifo_0_deqVld(cmdArbiter_io_fifo_0_deqVld),
    .io_fifo_0_empty(cmdArbiter_io_fifo_0_empty),
    .io_fifo_0_almostEmpty(cmdArbiter_io_fifo_0_almostEmpty),
    .io_fifo_1_deq_0_addr(cmdArbiter_io_fifo_1_deq_0_addr),
    .io_fifo_1_deq_0_isWr(cmdArbiter_io_fifo_1_deq_0_isWr),
    .io_fifo_1_deq_0_size(cmdArbiter_io_fifo_1_deq_0_size),
    .io_fifo_1_deqVld(cmdArbiter_io_fifo_1_deqVld),
    .io_fifo_1_empty(cmdArbiter_io_fifo_1_empty),
    .io_deq_0_addr(cmdArbiter_io_deq_0_addr),
    .io_deq_0_isWr(cmdArbiter_io_deq_0_isWr),
    .io_deq_0_size(cmdArbiter_io_deq_0_size),
    .io_deqVld(cmdArbiter_io_deqVld),
    .io_empty(cmdArbiter_io_empty),
    .io_tag(cmdArbiter_io_tag)
  );
  FIFOCore cmdFifos_0 (
    .clock(cmdFifos_0_clock),
    .reset(cmdFifos_0_reset),
    .io_deq_0_addr(cmdFifos_0_io_deq_0_addr),
    .io_deq_0_isWr(cmdFifos_0_io_deq_0_isWr),
    .io_deq_0_size(cmdFifos_0_io_deq_0_size),
    .io_deqVld(cmdFifos_0_io_deqVld),
    .io_empty(cmdFifos_0_io_empty),
    .io_almostEmpty(cmdFifos_0_io_almostEmpty)
  );
  FIFOCore cmdFifos_1 (
    .clock(cmdFifos_1_clock),
    .reset(cmdFifos_1_reset),
    .io_deq_0_addr(cmdFifos_1_io_deq_0_addr),
    .io_deq_0_isWr(cmdFifos_1_io_deq_0_isWr),
    .io_deq_0_size(cmdFifos_1_io_deq_0_size),
    .io_deqVld(cmdFifos_1_io_deqVld),
    .io_empty(cmdFifos_1_io_empty),
    .io_almostEmpty(cmdFifos_1_io_almostEmpty)
  );
  Counter_8 burstCounter (
    .clock(burstCounter_clock),
    .reset(burstCounter_reset),
    .io_max(burstCounter_io_max),
    .io_out(burstCounter_io_out),
    .io_enable(burstCounter_io_enable),
    .io_done(burstCounter_io_done)
  );
  Counter burstTagCounter (
    .clock(burstTagCounter_clock),
    .reset(burstTagCounter_reset),
    .io_max(burstTagCounter_io_max),
    .io_out(burstTagCounter_io_out),
    .io_next(burstTagCounter_io_next),
    .io_enable(burstTagCounter_io_enable),
    .io_done(burstTagCounter_io_done)
  );
  MuxN_3 rrespReadyMux (
    .io_ins_0(rrespReadyMux_io_ins_0),
    .io_out(rrespReadyMux_io_out)
  );
  MuxN_4 wdataMux (
    .io_ins_0_valid(wdataMux_io_ins_0_valid),
    .io_ins_0_bits_wdata_0(wdataMux_io_ins_0_bits_wdata_0),
    .io_ins_0_bits_wdata_1(wdataMux_io_ins_0_bits_wdata_1),
    .io_ins_0_bits_wdata_2(wdataMux_io_ins_0_bits_wdata_2),
    .io_ins_0_bits_wdata_3(wdataMux_io_ins_0_bits_wdata_3),
    .io_ins_0_bits_wdata_4(wdataMux_io_ins_0_bits_wdata_4),
    .io_ins_0_bits_wdata_5(wdataMux_io_ins_0_bits_wdata_5),
    .io_ins_0_bits_wdata_6(wdataMux_io_ins_0_bits_wdata_6),
    .io_ins_0_bits_wdata_7(wdataMux_io_ins_0_bits_wdata_7),
    .io_ins_0_bits_wdata_8(wdataMux_io_ins_0_bits_wdata_8),
    .io_ins_0_bits_wdata_9(wdataMux_io_ins_0_bits_wdata_9),
    .io_ins_0_bits_wdata_10(wdataMux_io_ins_0_bits_wdata_10),
    .io_ins_0_bits_wdata_11(wdataMux_io_ins_0_bits_wdata_11),
    .io_ins_0_bits_wdata_12(wdataMux_io_ins_0_bits_wdata_12),
    .io_ins_0_bits_wdata_13(wdataMux_io_ins_0_bits_wdata_13),
    .io_ins_0_bits_wdata_14(wdataMux_io_ins_0_bits_wdata_14),
    .io_ins_0_bits_wdata_15(wdataMux_io_ins_0_bits_wdata_15),
    .io_ins_0_bits_wlast(wdataMux_io_ins_0_bits_wlast),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wlast(wdataMux_io_out_bits_wlast)
  );
  MuxN_5 cmdDeqValidMux (
    .io_ins_0(cmdDeqValidMux_io_ins_0),
    .io_ins_1(cmdDeqValidMux_io_ins_1),
    .io_sel(cmdDeqValidMux_io_sel),
    .io_out(cmdDeqValidMux_io_out)
  );
  MuxN_6 dramCmdMux (
    .io_ins_0_valid(dramCmdMux_io_ins_0_valid),
    .io_ins_0_bits_addr(dramCmdMux_io_ins_0_bits_addr),
    .io_ins_0_bits_size(dramCmdMux_io_ins_0_bits_size),
    .io_ins_0_bits_isWr(dramCmdMux_io_ins_0_bits_isWr),
    .io_ins_0_bits_tag_uid(dramCmdMux_io_ins_0_bits_tag_uid),
    .io_ins_0_bits_tag_streamId(dramCmdMux_io_ins_0_bits_tag_streamId),
    .io_ins_1_valid(dramCmdMux_io_ins_1_valid),
    .io_ins_1_bits_addr(dramCmdMux_io_ins_1_bits_addr),
    .io_ins_1_bits_size(dramCmdMux_io_ins_1_bits_size),
    .io_ins_1_bits_isWr(dramCmdMux_io_ins_1_bits_isWr),
    .io_ins_1_bits_tag_uid(dramCmdMux_io_ins_1_bits_tag_uid),
    .io_ins_1_bits_tag_streamId(dramCmdMux_io_ins_1_bits_tag_streamId),
    .io_sel(dramCmdMux_io_sel),
    .io_out_valid(dramCmdMux_io_out_valid),
    .io_out_bits_addr(dramCmdMux_io_out_bits_addr),
    .io_out_bits_size(dramCmdMux_io_out_bits_size),
    .io_out_bits_isWr(dramCmdMux_io_out_bits_isWr),
    .io_out_bits_tag_uid(dramCmdMux_io_out_bits_tag_uid),
    .io_out_bits_tag_streamId(dramCmdMux_io_out_bits_tag_streamId)
  );
  FF_25 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_in(FF_io_in),
    .io_init(FF_io_init),
    .io_out(FF_io_out),
    .io_enable(FF_io_enable)
  );
  FF_26 FF_1 (
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_in(FF_1_io_in),
    .io_init(FF_1_io_init),
    .io_out(FF_1_io_out),
    .io_enable(FF_1_io_enable)
  );
  FF_23 FF_2 (
    .clock(FF_2_clock),
    .reset(FF_2_reset),
    .io_in(FF_2_io_in),
    .io_init(FF_2_io_init),
    .io_out(FF_2_io_out),
    .io_enable(FF_2_io_enable)
  );
  FF_2 FF_3 (
    .clock(FF_3_clock),
    .reset(FF_3_reset),
    .io_in(FF_3_io_in),
    .io_init(FF_3_io_init),
    .io_out(FF_3_io_out),
    .io_enable(FF_3_io_enable)
  );
  FF_26 FF_4 (
    .clock(FF_4_clock),
    .reset(FF_4_reset),
    .io_in(FF_4_io_in),
    .io_init(FF_4_io_init),
    .io_out(FF_4_io_out),
    .io_enable(FF_4_io_enable)
  );
  FF_30 FF_5 (
    .clock(FF_5_clock),
    .reset(FF_5_reset),
    .io_in(FF_5_io_in),
    .io_out(FF_5_io_out),
    .io_enable(FF_5_io_enable)
  );
  MuxN_3 wrespReadyMux (
    .io_ins_0(wrespReadyMux_io_ins_0),
    .io_out(wrespReadyMux_io_out)
  );
  MuxN_5 gatherLoadIssueMux (
    .io_ins_0(gatherLoadIssueMux_io_ins_0),
    .io_ins_1(gatherLoadIssueMux_io_ins_1),
    .io_sel(gatherLoadIssueMux_io_sel),
    .io_out(gatherLoadIssueMux_io_out)
  );
  Counter_8 gatherLoadIssue (
    .clock(gatherLoadIssue_clock),
    .reset(gatherLoadIssue_reset),
    .io_max(gatherLoadIssue_io_max),
    .io_out(gatherLoadIssue_io_out),
    .io_enable(gatherLoadIssue_io_enable),
    .io_done(gatherLoadIssue_io_done)
  );
  MuxN_5 gatherLoadSkipMux (
    .io_ins_0(gatherLoadSkipMux_io_ins_0),
    .io_ins_1(gatherLoadSkipMux_io_ins_1),
    .io_sel(gatherLoadSkipMux_io_sel),
    .io_out(gatherLoadSkipMux_io_out)
  );
  Counter_8 gatherLoadSkip (
    .clock(gatherLoadSkip_clock),
    .reset(gatherLoadSkip_reset),
    .io_max(gatherLoadSkip_io_max),
    .io_out(gatherLoadSkip_io_out),
    .io_enable(gatherLoadSkip_io_enable),
    .io_done(gatherLoadSkip_io_done)
  );
  MuxN_5 scatterLoadIssueMux (
    .io_ins_0(scatterLoadIssueMux_io_ins_0),
    .io_ins_1(scatterLoadIssueMux_io_ins_1),
    .io_sel(scatterLoadIssueMux_io_sel),
    .io_out(scatterLoadIssueMux_io_out)
  );
  Counter_8 scatterLoadIssue (
    .clock(scatterLoadIssue_clock),
    .reset(scatterLoadIssue_reset),
    .io_max(scatterLoadIssue_io_max),
    .io_out(scatterLoadIssue_io_out),
    .io_enable(scatterLoadIssue_io_enable),
    .io_done(scatterLoadIssue_io_done)
  );
  MuxN_5 scatterLoadSkipMux (
    .io_ins_0(scatterLoadSkipMux_io_ins_0),
    .io_ins_1(scatterLoadSkipMux_io_ins_1),
    .io_sel(scatterLoadSkipMux_io_sel),
    .io_out(scatterLoadSkipMux_io_out)
  );
  Counter_8 scatterLoadSkip (
    .clock(scatterLoadSkip_clock),
    .reset(scatterLoadSkip_reset),
    .io_max(scatterLoadSkip_io_max),
    .io_out(scatterLoadSkip_io_out),
    .io_enable(scatterLoadSkip_io_enable),
    .io_done(scatterLoadSkip_io_done)
  );
  MuxN_5 scatterStoreIssueMux (
    .io_ins_0(scatterStoreIssueMux_io_ins_0),
    .io_ins_1(scatterStoreIssueMux_io_ins_1),
    .io_sel(scatterStoreIssueMux_io_sel),
    .io_out(scatterStoreIssueMux_io_out)
  );
  Counter_8 scatterStoreIssue (
    .clock(scatterStoreIssue_clock),
    .reset(scatterStoreIssue_reset),
    .io_max(scatterStoreIssue_io_max),
    .io_out(scatterStoreIssue_io_out),
    .io_enable(scatterStoreIssue_io_enable),
    .io_done(scatterStoreIssue_io_done)
  );
  MuxN_5 scatterStoreSkipMux (
    .io_ins_0(scatterStoreSkipMux_io_ins_0),
    .io_ins_1(scatterStoreSkipMux_io_ins_1),
    .io_sel(scatterStoreSkipMux_io_sel),
    .io_out(scatterStoreSkipMux_io_out)
  );
  Counter_8 scatterStoreSkip (
    .clock(scatterStoreSkip_clock),
    .reset(scatterStoreSkip_reset),
    .io_max(scatterStoreSkip_io_max),
    .io_out(scatterStoreSkip_io_out),
    .io_enable(scatterStoreSkip_io_enable),
    .io_done(scatterStoreSkip_io_done)
  );
  FIFOWidthConvert denseLoadBuffers_0 (
    .clock(denseLoadBuffers_0_clock),
    .reset(denseLoadBuffers_0_reset),
    .io_enq_0(denseLoadBuffers_0_io_enq_0),
    .io_enq_1(denseLoadBuffers_0_io_enq_1),
    .io_enq_2(denseLoadBuffers_0_io_enq_2),
    .io_enq_3(denseLoadBuffers_0_io_enq_3),
    .io_enq_4(denseLoadBuffers_0_io_enq_4),
    .io_enq_5(denseLoadBuffers_0_io_enq_5),
    .io_enq_6(denseLoadBuffers_0_io_enq_6),
    .io_enq_7(denseLoadBuffers_0_io_enq_7),
    .io_enq_8(denseLoadBuffers_0_io_enq_8),
    .io_enq_9(denseLoadBuffers_0_io_enq_9),
    .io_enq_10(denseLoadBuffers_0_io_enq_10),
    .io_enq_11(denseLoadBuffers_0_io_enq_11),
    .io_enq_12(denseLoadBuffers_0_io_enq_12),
    .io_enq_13(denseLoadBuffers_0_io_enq_13),
    .io_enq_14(denseLoadBuffers_0_io_enq_14),
    .io_enq_15(denseLoadBuffers_0_io_enq_15),
    .io_enqVld(denseLoadBuffers_0_io_enqVld),
    .io_deq_0(denseLoadBuffers_0_io_deq_0),
    .io_deq_1(denseLoadBuffers_0_io_deq_1),
    .io_deq_2(denseLoadBuffers_0_io_deq_2),
    .io_deq_3(denseLoadBuffers_0_io_deq_3),
    .io_deq_4(denseLoadBuffers_0_io_deq_4),
    .io_deq_5(denseLoadBuffers_0_io_deq_5),
    .io_deq_6(denseLoadBuffers_0_io_deq_6),
    .io_deq_7(denseLoadBuffers_0_io_deq_7),
    .io_deq_8(denseLoadBuffers_0_io_deq_8),
    .io_deq_9(denseLoadBuffers_0_io_deq_9),
    .io_deq_10(denseLoadBuffers_0_io_deq_10),
    .io_deq_11(denseLoadBuffers_0_io_deq_11),
    .io_deq_12(denseLoadBuffers_0_io_deq_12),
    .io_deq_13(denseLoadBuffers_0_io_deq_13),
    .io_deq_14(denseLoadBuffers_0_io_deq_14),
    .io_deq_15(denseLoadBuffers_0_io_deq_15),
    .io_deqVld(denseLoadBuffers_0_io_deqVld),
    .io_full(denseLoadBuffers_0_io_full),
    .io_empty(denseLoadBuffers_0_io_empty),
    .io_almostEmpty(denseLoadBuffers_0_io_almostEmpty),
    .io_almostFull(denseLoadBuffers_0_io_almostFull)
  );
  Counter_8 Counter (
    .clock(Counter_clock),
    .reset(Counter_reset),
    .io_max(Counter_io_max),
    .io_out(Counter_io_out),
    .io_enable(Counter_io_enable),
    .io_done(Counter_io_done)
  );
  Counter_8 Counter_1 (
    .clock(Counter_1_clock),
    .reset(Counter_1_reset),
    .io_max(Counter_1_io_max),
    .io_out(Counter_1_io_out),
    .io_enable(Counter_1_io_enable),
    .io_done(Counter_1_io_done)
  );
  SRFF_sp SRFF_sp (
    .clock(SRFF_sp_clock),
    .reset(SRFF_sp_reset),
    .io_input_set(SRFF_sp_io_input_set),
    .io_input_reset(SRFF_sp_io_input_reset),
    .io_input_asyn_reset(SRFF_sp_io_input_asyn_reset),
    .io_output_data(SRFF_sp_io_output_data)
  );
  SRFF_sp SRFF_sp_1 (
    .clock(SRFF_sp_1_clock),
    .reset(SRFF_sp_1_reset),
    .io_input_set(SRFF_sp_1_io_input_set),
    .io_input_reset(SRFF_sp_1_io_input_reset),
    .io_input_asyn_reset(SRFF_sp_1_io_input_asyn_reset),
    .io_output_data(SRFF_sp_1_io_output_data)
  );
  FF_49 FF_6 (
    .clock(FF_6_clock),
    .reset(FF_6_reset),
    .io_in(FF_6_io_in),
    .io_init(FF_6_io_init),
    .io_out(FF_6_io_out),
    .io_enable(FF_6_io_enable)
  );
  FF_49 FF_7 (
    .clock(FF_7_clock),
    .reset(FF_7_reset),
    .io_in(FF_7_io_in),
    .io_init(FF_7_io_init),
    .io_out(FF_7_io_out),
    .io_enable(FF_7_io_enable)
  );
  FIFOWidthConvert denseStoreBuffers_0 (
    .clock(denseStoreBuffers_0_clock),
    .reset(denseStoreBuffers_0_reset),
    .io_enq_0(denseStoreBuffers_0_io_enq_0),
    .io_enq_1(denseStoreBuffers_0_io_enq_1),
    .io_enq_2(denseStoreBuffers_0_io_enq_2),
    .io_enq_3(denseStoreBuffers_0_io_enq_3),
    .io_enq_4(denseStoreBuffers_0_io_enq_4),
    .io_enq_5(denseStoreBuffers_0_io_enq_5),
    .io_enq_6(denseStoreBuffers_0_io_enq_6),
    .io_enq_7(denseStoreBuffers_0_io_enq_7),
    .io_enq_8(denseStoreBuffers_0_io_enq_8),
    .io_enq_9(denseStoreBuffers_0_io_enq_9),
    .io_enq_10(denseStoreBuffers_0_io_enq_10),
    .io_enq_11(denseStoreBuffers_0_io_enq_11),
    .io_enq_12(denseStoreBuffers_0_io_enq_12),
    .io_enq_13(denseStoreBuffers_0_io_enq_13),
    .io_enq_14(denseStoreBuffers_0_io_enq_14),
    .io_enq_15(denseStoreBuffers_0_io_enq_15),
    .io_enqVld(denseStoreBuffers_0_io_enqVld),
    .io_deq_0(denseStoreBuffers_0_io_deq_0),
    .io_deq_1(denseStoreBuffers_0_io_deq_1),
    .io_deq_2(denseStoreBuffers_0_io_deq_2),
    .io_deq_3(denseStoreBuffers_0_io_deq_3),
    .io_deq_4(denseStoreBuffers_0_io_deq_4),
    .io_deq_5(denseStoreBuffers_0_io_deq_5),
    .io_deq_6(denseStoreBuffers_0_io_deq_6),
    .io_deq_7(denseStoreBuffers_0_io_deq_7),
    .io_deq_8(denseStoreBuffers_0_io_deq_8),
    .io_deq_9(denseStoreBuffers_0_io_deq_9),
    .io_deq_10(denseStoreBuffers_0_io_deq_10),
    .io_deq_11(denseStoreBuffers_0_io_deq_11),
    .io_deq_12(denseStoreBuffers_0_io_deq_12),
    .io_deq_13(denseStoreBuffers_0_io_deq_13),
    .io_deq_14(denseStoreBuffers_0_io_deq_14),
    .io_deq_15(denseStoreBuffers_0_io_deq_15),
    .io_deqVld(denseStoreBuffers_0_io_deqVld),
    .io_full(denseStoreBuffers_0_io_full),
    .io_empty(denseStoreBuffers_0_io_empty),
    .io_almostEmpty(denseStoreBuffers_0_io_almostEmpty),
    .io_almostFull(denseStoreBuffers_0_io_almostFull)
  );
  FIFOCounter FIFOCounter (
    .clock(FIFOCounter_clock),
    .reset(FIFOCounter_reset),
    .io_enqVld(FIFOCounter_io_enqVld),
    .io_full(FIFOCounter_io_full)
  );
  Counter_8 Counter_2 (
    .clock(Counter_2_clock),
    .reset(Counter_2_reset),
    .io_max(Counter_2_io_max),
    .io_out(Counter_2_io_out),
    .io_enable(Counter_2_io_enable),
    .io_done(Counter_2_io_done)
  );
  FFType dramReadyFF (
    .clock(dramReadyFF_clock),
    .reset(dramReadyFF_reset),
    .io_in(dramReadyFF_io_in),
    .io_init(dramReadyFF_io_init),
    .io_out(dramReadyFF_io_out),
    .io_enable(dramReadyFF_io_enable)
  );
  Counter_8 cycleCount (
    .clock(cycleCount_clock),
    .reset(cycleCount_reset),
    .io_max(cycleCount_io_max),
    .io_out(cycleCount_io_out),
    .io_enable(cycleCount_io_enable),
    .io_done(cycleCount_io_done)
  );
  Counter_8 rdataEnqCount (
    .clock(rdataEnqCount_clock),
    .reset(rdataEnqCount_reset),
    .io_max(rdataEnqCount_io_max),
    .io_out(rdataEnqCount_io_out),
    .io_enable(rdataEnqCount_io_enable),
    .io_done(rdataEnqCount_io_done)
  );
  Counter_8 wdataCount (
    .clock(wdataCount_clock),
    .reset(wdataCount_reset),
    .io_max(wdataCount_io_max),
    .io_out(wdataCount_io_out),
    .io_enable(wdataCount_io_enable),
    .io_done(wdataCount_io_done)
  );
  FF_23 FF_8 (
    .clock(FF_8_clock),
    .reset(FF_8_reset),
    .io_in(FF_8_io_in),
    .io_init(FF_8_io_init),
    .io_out(FF_8_io_out),
    .io_enable(FF_8_io_enable)
  );
  FF_23 FF_9 (
    .clock(FF_9_clock),
    .reset(FF_9_reset),
    .io_in(FF_9_io_in),
    .io_init(FF_9_io_init),
    .io_out(FF_9_io_out),
    .io_enable(FF_9_io_enable)
  );
  FF_23 FF_10 (
    .clock(FF_10_clock),
    .reset(FF_10_reset),
    .io_in(FF_10_io_in),
    .io_init(FF_10_io_init),
    .io_out(FF_10_io_out),
    .io_enable(FF_10_io_enable)
  );
  FF_23 FF_11 (
    .clock(FF_11_clock),
    .reset(FF_11_reset),
    .io_in(FF_11_io_in),
    .io_init(FF_11_io_init),
    .io_out(FF_11_io_out),
    .io_enable(FF_11_io_enable)
  );
  FF_23 FF_12 (
    .clock(FF_12_clock),
    .reset(FF_12_reset),
    .io_in(FF_12_io_in),
    .io_init(FF_12_io_init),
    .io_out(FF_12_io_out),
    .io_enable(FF_12_io_enable)
  );
  FF_23 FF_13 (
    .clock(FF_13_clock),
    .reset(FF_13_reset),
    .io_in(FF_13_io_in),
    .io_init(FF_13_io_init),
    .io_out(FF_13_io_out),
    .io_enable(FF_13_io_enable)
  );
  FF_23 FF_14 (
    .clock(FF_14_clock),
    .reset(FF_14_reset),
    .io_in(FF_14_io_in),
    .io_init(FF_14_io_init),
    .io_out(FF_14_io_out),
    .io_enable(FF_14_io_enable)
  );
  FF_23 FF_15 (
    .clock(FF_15_clock),
    .reset(FF_15_reset),
    .io_in(FF_15_io_in),
    .io_init(FF_15_io_init),
    .io_out(FF_15_io_out),
    .io_enable(FF_15_io_enable)
  );
  FF_23 FF_16 (
    .clock(FF_16_clock),
    .reset(FF_16_reset),
    .io_in(FF_16_io_in),
    .io_init(FF_16_io_init),
    .io_out(FF_16_io_out),
    .io_enable(FF_16_io_enable)
  );
  FF_23 FF_17 (
    .clock(FF_17_clock),
    .reset(FF_17_reset),
    .io_in(FF_17_io_in),
    .io_init(FF_17_io_init),
    .io_out(FF_17_io_out),
    .io_enable(FF_17_io_enable)
  );
  FF_23 FF_18 (
    .clock(FF_18_clock),
    .reset(FF_18_reset),
    .io_in(FF_18_io_in),
    .io_init(FF_18_io_init),
    .io_out(FF_18_io_out),
    .io_enable(FF_18_io_enable)
  );
  FF_23 FF_19 (
    .clock(FF_19_clock),
    .reset(FF_19_reset),
    .io_in(FF_19_io_in),
    .io_init(FF_19_io_init),
    .io_out(FF_19_io_out),
    .io_enable(FF_19_io_enable)
  );
  FF_23 FF_20 (
    .clock(FF_20_clock),
    .reset(FF_20_reset),
    .io_in(FF_20_io_in),
    .io_init(FF_20_io_init),
    .io_out(FF_20_io_out),
    .io_enable(FF_20_io_enable)
  );
  FF_23 FF_21 (
    .clock(FF_21_clock),
    .reset(FF_21_reset),
    .io_in(FF_21_io_in),
    .io_init(FF_21_io_init),
    .io_out(FF_21_io_out),
    .io_enable(FF_21_io_enable)
  );
  FF_23 FF_22 (
    .clock(FF_22_clock),
    .reset(FF_22_reset),
    .io_in(FF_22_io_in),
    .io_init(FF_22_io_init),
    .io_out(FF_22_io_out),
    .io_enable(FF_22_io_enable)
  );
  FF_23 FF_23 (
    .clock(FF_23_clock),
    .reset(FF_23_reset),
    .io_in(FF_23_io_in),
    .io_init(FF_23_io_init),
    .io_out(FF_23_io_out),
    .io_enable(FF_23_io_enable)
  );
  FF_23 FF_24 (
    .clock(FF_24_clock),
    .reset(FF_24_reset),
    .io_in(FF_24_io_in),
    .io_init(FF_24_io_init),
    .io_out(FF_24_io_out),
    .io_enable(FF_24_io_enable)
  );
  FF_23 FF_25 (
    .clock(FF_25_clock),
    .reset(FF_25_reset),
    .io_in(FF_25_io_in),
    .io_init(FF_25_io_init),
    .io_out(FF_25_io_out),
    .io_enable(FF_25_io_enable)
  );
  FF_23 FF_26 (
    .clock(FF_26_clock),
    .reset(FF_26_reset),
    .io_in(FF_26_io_in),
    .io_init(FF_26_io_init),
    .io_out(FF_26_io_out),
    .io_enable(FF_26_io_enable)
  );
  FF_23 FF_27 (
    .clock(FF_27_clock),
    .reset(FF_27_reset),
    .io_in(FF_27_io_in),
    .io_init(FF_27_io_init),
    .io_out(FF_27_io_out),
    .io_enable(FF_27_io_enable)
  );
  FF_23 FF_28 (
    .clock(FF_28_clock),
    .reset(FF_28_reset),
    .io_in(FF_28_io_in),
    .io_init(FF_28_io_init),
    .io_out(FF_28_io_out),
    .io_enable(FF_28_io_enable)
  );
  FF_23 FF_29 (
    .clock(FF_29_clock),
    .reset(FF_29_reset),
    .io_in(FF_29_io_in),
    .io_init(FF_29_io_init),
    .io_out(FF_29_io_out),
    .io_enable(FF_29_io_enable)
  );
  FF_23 FF_30 (
    .clock(FF_30_clock),
    .reset(FF_30_reset),
    .io_in(FF_30_io_in),
    .io_init(FF_30_io_init),
    .io_out(FF_30_io_out),
    .io_enable(FF_30_io_enable)
  );
  FF_23 FF_31 (
    .clock(FF_31_clock),
    .reset(FF_31_reset),
    .io_in(FF_31_io_in),
    .io_init(FF_31_io_init),
    .io_out(FF_31_io_out),
    .io_enable(FF_31_io_enable)
  );
  FF_23 FF_32 (
    .clock(FF_32_clock),
    .reset(FF_32_reset),
    .io_in(FF_32_io_in),
    .io_init(FF_32_io_init),
    .io_out(FF_32_io_out),
    .io_enable(FF_32_io_enable)
  );
  FF_23 FF_33 (
    .clock(FF_33_clock),
    .reset(FF_33_reset),
    .io_in(FF_33_io_in),
    .io_init(FF_33_io_init),
    .io_out(FF_33_io_out),
    .io_enable(FF_33_io_enable)
  );
  FF_23 FF_34 (
    .clock(FF_34_clock),
    .reset(FF_34_reset),
    .io_in(FF_34_io_in),
    .io_init(FF_34_io_init),
    .io_out(FF_34_io_out),
    .io_enable(FF_34_io_enable)
  );
  FF_23 FF_35 (
    .clock(FF_35_clock),
    .reset(FF_35_reset),
    .io_in(FF_35_io_in),
    .io_init(FF_35_io_init),
    .io_out(FF_35_io_out),
    .io_enable(FF_35_io_enable)
  );
  FF_23 FF_36 (
    .clock(FF_36_clock),
    .reset(FF_36_reset),
    .io_in(FF_36_io_in),
    .io_init(FF_36_io_init),
    .io_out(FF_36_io_out),
    .io_enable(FF_36_io_enable)
  );
  FF_23 FF_37 (
    .clock(FF_37_clock),
    .reset(FF_37_reset),
    .io_in(FF_37_io_in),
    .io_init(FF_37_io_init),
    .io_out(FF_37_io_out),
    .io_enable(FF_37_io_enable)
  );
  FF_23 FF_38 (
    .clock(FF_38_clock),
    .reset(FF_38_reset),
    .io_in(FF_38_io_in),
    .io_init(FF_38_io_init),
    .io_out(FF_38_io_out),
    .io_enable(FF_38_io_enable)
  );
  FF_23 FF_39 (
    .clock(FF_39_clock),
    .reset(FF_39_reset),
    .io_in(FF_39_io_in),
    .io_init(FF_39_io_init),
    .io_out(FF_39_io_out),
    .io_enable(FF_39_io_enable)
  );
  FF_23 FF_40 (
    .clock(FF_40_clock),
    .reset(FF_40_reset),
    .io_in(FF_40_io_in),
    .io_init(FF_40_io_init),
    .io_out(FF_40_io_out),
    .io_enable(FF_40_io_enable)
  );
  FF_23 FF_41 (
    .clock(FF_41_clock),
    .reset(FF_41_reset),
    .io_in(FF_41_io_in),
    .io_init(FF_41_io_init),
    .io_out(FF_41_io_out),
    .io_enable(FF_41_io_enable)
  );
  FF_23 FF_42 (
    .clock(FF_42_clock),
    .reset(FF_42_reset),
    .io_in(FF_42_io_in),
    .io_init(FF_42_io_init),
    .io_out(FF_42_io_out),
    .io_enable(FF_42_io_enable)
  );
  FF_23 FF_43 (
    .clock(FF_43_clock),
    .reset(FF_43_reset),
    .io_in(FF_43_io_in),
    .io_init(FF_43_io_init),
    .io_out(FF_43_io_out),
    .io_enable(FF_43_io_enable)
  );
  FF_23 FF_44 (
    .clock(FF_44_clock),
    .reset(FF_44_reset),
    .io_in(FF_44_io_in),
    .io_init(FF_44_io_init),
    .io_out(FF_44_io_out),
    .io_enable(FF_44_io_enable)
  );
  FF_23 FF_45 (
    .clock(FF_45_clock),
    .reset(FF_45_reset),
    .io_in(FF_45_io_in),
    .io_init(FF_45_io_init),
    .io_out(FF_45_io_out),
    .io_enable(FF_45_io_enable)
  );
  FF_23 FF_46 (
    .clock(FF_46_clock),
    .reset(FF_46_reset),
    .io_in(FF_46_io_in),
    .io_init(FF_46_io_init),
    .io_out(FF_46_io_out),
    .io_enable(FF_46_io_enable)
  );
  FF_23 FF_47 (
    .clock(FF_47_clock),
    .reset(FF_47_reset),
    .io_in(FF_47_io_in),
    .io_init(FF_47_io_init),
    .io_out(FF_47_io_out),
    .io_enable(FF_47_io_enable)
  );
  FF_23 FF_48 (
    .clock(FF_48_clock),
    .reset(FF_48_reset),
    .io_in(FF_48_io_in),
    .io_init(FF_48_io_init),
    .io_out(FF_48_io_out),
    .io_enable(FF_48_io_enable)
  );
  FF_23 FF_49 (
    .clock(FF_49_clock),
    .reset(FF_49_reset),
    .io_in(FF_49_io_in),
    .io_init(FF_49_io_init),
    .io_out(FF_49_io_out),
    .io_enable(FF_49_io_enable)
  );
  FF_23 FF_50 (
    .clock(FF_50_clock),
    .reset(FF_50_reset),
    .io_in(FF_50_io_in),
    .io_init(FF_50_io_init),
    .io_out(FF_50_io_out),
    .io_enable(FF_50_io_enable)
  );
  FF_23 FF_51 (
    .clock(FF_51_clock),
    .reset(FF_51_reset),
    .io_in(FF_51_io_in),
    .io_init(FF_51_io_init),
    .io_out(FF_51_io_out),
    .io_enable(FF_51_io_enable)
  );
  FF_23 FF_52 (
    .clock(FF_52_clock),
    .reset(FF_52_reset),
    .io_in(FF_52_io_in),
    .io_init(FF_52_io_init),
    .io_out(FF_52_io_out),
    .io_enable(FF_52_io_enable)
  );
  FF_23 FF_53 (
    .clock(FF_53_clock),
    .reset(FF_53_reset),
    .io_in(FF_53_io_in),
    .io_init(FF_53_io_init),
    .io_out(FF_53_io_out),
    .io_enable(FF_53_io_enable)
  );
  FF_23 FF_54 (
    .clock(FF_54_clock),
    .reset(FF_54_reset),
    .io_in(FF_54_io_in),
    .io_init(FF_54_io_init),
    .io_out(FF_54_io_out),
    .io_enable(FF_54_io_enable)
  );
  FF_23 FF_55 (
    .clock(FF_55_clock),
    .reset(FF_55_reset),
    .io_in(FF_55_io_in),
    .io_init(FF_55_io_init),
    .io_out(FF_55_io_out),
    .io_enable(FF_55_io_enable)
  );
  FF_49 FF_56 (
    .clock(FF_56_clock),
    .reset(FF_56_reset),
    .io_in(FF_56_io_in),
    .io_init(FF_56_io_init),
    .io_out(FF_56_io_out),
    .io_enable(FF_56_io_enable)
  );
  FF_23 FF_57 (
    .clock(FF_57_clock),
    .reset(FF_57_reset),
    .io_in(FF_57_io_in),
    .io_init(FF_57_io_init),
    .io_out(FF_57_io_out),
    .io_enable(FF_57_io_enable)
  );
  FF_23 FF_58 (
    .clock(FF_58_clock),
    .reset(FF_58_reset),
    .io_in(FF_58_io_in),
    .io_init(FF_58_io_init),
    .io_out(FF_58_io_out),
    .io_enable(FF_58_io_enable)
  );
  FF_23 FF_59 (
    .clock(FF_59_clock),
    .reset(FF_59_reset),
    .io_in(FF_59_io_in),
    .io_init(FF_59_io_init),
    .io_out(FF_59_io_out),
    .io_enable(FF_59_io_enable)
  );
  FF_23 FF_60 (
    .clock(FF_60_clock),
    .reset(FF_60_reset),
    .io_in(FF_60_io_in),
    .io_init(FF_60_io_init),
    .io_out(FF_60_io_out),
    .io_enable(FF_60_io_enable)
  );
  FF_23 FF_61 (
    .clock(FF_61_clock),
    .reset(FF_61_reset),
    .io_in(FF_61_io_in),
    .io_init(FF_61_io_init),
    .io_out(FF_61_io_out),
    .io_enable(FF_61_io_enable)
  );
  FF_23 FF_62 (
    .clock(FF_62_clock),
    .reset(FF_62_reset),
    .io_in(FF_62_io_in),
    .io_init(FF_62_io_init),
    .io_out(FF_62_io_out),
    .io_enable(FF_62_io_enable)
  );
  FF_23 FF_63 (
    .clock(FF_63_clock),
    .reset(FF_63_reset),
    .io_in(FF_63_io_in),
    .io_init(FF_63_io_init),
    .io_out(FF_63_io_out),
    .io_enable(FF_63_io_enable)
  );
  FF_23 FF_64 (
    .clock(FF_64_clock),
    .reset(FF_64_reset),
    .io_in(FF_64_io_in),
    .io_init(FF_64_io_init),
    .io_out(FF_64_io_out),
    .io_enable(FF_64_io_enable)
  );
  FF_23 FF_65 (
    .clock(FF_65_clock),
    .reset(FF_65_reset),
    .io_in(FF_65_io_in),
    .io_init(FF_65_io_init),
    .io_out(FF_65_io_out),
    .io_enable(FF_65_io_enable)
  );
  FF_23 FF_66 (
    .clock(FF_66_clock),
    .reset(FF_66_reset),
    .io_in(FF_66_io_in),
    .io_init(FF_66_io_init),
    .io_out(FF_66_io_out),
    .io_enable(FF_66_io_enable)
  );
  FF_23 FF_67 (
    .clock(FF_67_clock),
    .reset(FF_67_reset),
    .io_in(FF_67_io_in),
    .io_init(FF_67_io_init),
    .io_out(FF_67_io_out),
    .io_enable(FF_67_io_enable)
  );
  FF_23 FF_68 (
    .clock(FF_68_clock),
    .reset(FF_68_reset),
    .io_in(FF_68_io_in),
    .io_init(FF_68_io_init),
    .io_out(FF_68_io_out),
    .io_enable(FF_68_io_enable)
  );
  FF_23 FF_69 (
    .clock(FF_69_clock),
    .reset(FF_69_reset),
    .io_in(FF_69_io_in),
    .io_init(FF_69_io_init),
    .io_out(FF_69_io_out),
    .io_enable(FF_69_io_enable)
  );
  FF_23 FF_70 (
    .clock(FF_70_clock),
    .reset(FF_70_reset),
    .io_in(FF_70_io_in),
    .io_init(FF_70_io_init),
    .io_out(FF_70_io_out),
    .io_enable(FF_70_io_enable)
  );
  FF_23 FF_71 (
    .clock(FF_71_clock),
    .reset(FF_71_reset),
    .io_in(FF_71_io_in),
    .io_init(FF_71_io_init),
    .io_out(FF_71_io_out),
    .io_enable(FF_71_io_enable)
  );
  FF_23 FF_72 (
    .clock(FF_72_clock),
    .reset(FF_72_reset),
    .io_in(FF_72_io_in),
    .io_init(FF_72_io_init),
    .io_out(FF_72_io_out),
    .io_enable(FF_72_io_enable)
  );
  FF_49 FF_73 (
    .clock(FF_73_clock),
    .reset(FF_73_reset),
    .io_in(FF_73_io_in),
    .io_init(FF_73_io_init),
    .io_out(FF_73_io_out),
    .io_enable(FF_73_io_enable)
  );
  Counter_8 Counter_3 (
    .clock(Counter_3_clock),
    .reset(Counter_3_reset),
    .io_max(Counter_3_io_max),
    .io_out(Counter_3_io_out),
    .io_enable(Counter_3_io_enable),
    .io_done(Counter_3_io_done)
  );
  Counter_8 Counter_4 (
    .clock(Counter_4_clock),
    .reset(Counter_4_reset),
    .io_max(Counter_4_io_max),
    .io_out(Counter_4_io_out),
    .io_enable(Counter_4_io_enable),
    .io_done(Counter_4_io_done)
  );
  Counter_8 Counter_5 (
    .clock(Counter_5_clock),
    .reset(Counter_5_reset),
    .io_max(Counter_5_io_max),
    .io_out(Counter_5_io_out),
    .io_enable(Counter_5_io_enable),
    .io_done(Counter_5_io_done)
  );
  Counter_8 Counter_6 (
    .clock(Counter_6_clock),
    .reset(Counter_6_reset),
    .io_max(Counter_6_io_max),
    .io_out(Counter_6_io_out),
    .io_enable(Counter_6_io_enable),
    .io_done(Counter_6_io_done)
  );
  Counter_8 Counter_7 (
    .clock(Counter_7_clock),
    .reset(Counter_7_reset),
    .io_max(Counter_7_io_max),
    .io_out(Counter_7_io_out),
    .io_enable(Counter_7_io_enable),
    .io_done(Counter_7_io_done)
  );
  Counter_8 Counter_8 (
    .clock(Counter_8_clock),
    .reset(Counter_8_reset),
    .io_max(Counter_8_io_max),
    .io_out(Counter_8_io_out),
    .io_enable(Counter_8_io_enable),
    .io_done(Counter_8_io_done)
  );
  Counter_8 Counter_9 (
    .clock(Counter_9_clock),
    .reset(Counter_9_reset),
    .io_max(Counter_9_io_max),
    .io_out(Counter_9_io_out),
    .io_enable(Counter_9_io_enable),
    .io_done(Counter_9_io_done)
  );
  Counter_8 Counter_10 (
    .clock(Counter_10_clock),
    .reset(Counter_10_reset),
    .io_max(Counter_10_io_max),
    .io_out(Counter_10_io_out),
    .io_enable(Counter_10_io_enable),
    .io_done(Counter_10_io_done)
  );
  Counter_8 Counter_11 (
    .clock(Counter_11_clock),
    .reset(Counter_11_reset),
    .io_max(Counter_11_io_max),
    .io_out(Counter_11_io_out),
    .io_enable(Counter_11_io_enable),
    .io_done(Counter_11_io_done)
  );
  Counter_8 Counter_12 (
    .clock(Counter_12_clock),
    .reset(Counter_12_reset),
    .io_max(Counter_12_io_max),
    .io_out(Counter_12_io_out),
    .io_enable(Counter_12_io_enable),
    .io_done(Counter_12_io_done)
  );
  Counter_8 Counter_13 (
    .clock(Counter_13_clock),
    .reset(Counter_13_reset),
    .io_max(Counter_13_io_max),
    .io_out(Counter_13_io_out),
    .io_enable(Counter_13_io_enable),
    .io_done(Counter_13_io_done)
  );
  Counter_8 Counter_14 (
    .clock(Counter_14_clock),
    .reset(Counter_14_reset),
    .io_max(Counter_14_io_max),
    .io_out(Counter_14_io_out),
    .io_enable(Counter_14_io_enable),
    .io_done(Counter_14_io_done)
  );
  Counter_8 Counter_15 (
    .clock(Counter_15_clock),
    .reset(Counter_15_reset),
    .io_max(Counter_15_io_max),
    .io_out(Counter_15_io_out),
    .io_enable(Counter_15_io_enable),
    .io_done(Counter_15_io_done)
  );
  Counter_8 Counter_16 (
    .clock(Counter_16_clock),
    .reset(Counter_16_reset),
    .io_max(Counter_16_io_max),
    .io_out(Counter_16_io_out),
    .io_enable(Counter_16_io_enable),
    .io_done(Counter_16_io_done)
  );
  Counter_8 Counter_17 (
    .clock(Counter_17_clock),
    .reset(Counter_17_reset),
    .io_max(Counter_17_io_max),
    .io_out(Counter_17_io_out),
    .io_enable(Counter_17_io_enable),
    .io_done(Counter_17_io_done)
  );
  Counter_8 Counter_18 (
    .clock(Counter_18_clock),
    .reset(Counter_18_reset),
    .io_max(Counter_18_io_max),
    .io_out(Counter_18_io_out),
    .io_enable(Counter_18_io_enable),
    .io_done(Counter_18_io_done)
  );
  Counter_8 Counter_19 (
    .clock(Counter_19_clock),
    .reset(Counter_19_reset),
    .io_max(Counter_19_io_max),
    .io_out(Counter_19_io_out),
    .io_enable(Counter_19_io_enable),
    .io_done(Counter_19_io_done)
  );
  Counter_8 Counter_20 (
    .clock(Counter_20_clock),
    .reset(Counter_20_reset),
    .io_max(Counter_20_io_max),
    .io_out(Counter_20_io_out),
    .io_enable(Counter_20_io_enable),
    .io_done(Counter_20_io_done)
  );
  Counter_8 Counter_21 (
    .clock(Counter_21_clock),
    .reset(Counter_21_reset),
    .io_max(Counter_21_io_max),
    .io_out(Counter_21_io_out),
    .io_enable(Counter_21_io_enable),
    .io_done(Counter_21_io_done)
  );
  Counter_8 Counter_22 (
    .clock(Counter_22_clock),
    .reset(Counter_22_reset),
    .io_max(Counter_22_io_max),
    .io_out(Counter_22_io_out),
    .io_enable(Counter_22_io_enable),
    .io_done(Counter_22_io_done)
  );
  Counter_8 Counter_23 (
    .clock(Counter_23_clock),
    .reset(Counter_23_reset),
    .io_max(Counter_23_io_max),
    .io_out(Counter_23_io_out),
    .io_enable(Counter_23_io_enable),
    .io_done(Counter_23_io_done)
  );
  Counter_8 Counter_24 (
    .clock(Counter_24_clock),
    .reset(Counter_24_reset),
    .io_max(Counter_24_io_max),
    .io_out(Counter_24_io_out),
    .io_enable(Counter_24_io_enable),
    .io_done(Counter_24_io_done)
  );
  Counter_8 Counter_25 (
    .clock(Counter_25_clock),
    .reset(Counter_25_reset),
    .io_max(Counter_25_io_max),
    .io_out(Counter_25_io_out),
    .io_enable(Counter_25_io_enable),
    .io_done(Counter_25_io_done)
  );
  Counter_8 Counter_26 (
    .clock(Counter_26_clock),
    .reset(Counter_26_reset),
    .io_max(Counter_26_io_max),
    .io_out(Counter_26_io_out),
    .io_enable(Counter_26_io_enable),
    .io_done(Counter_26_io_done)
  );
  Counter_8 Counter_27 (
    .clock(Counter_27_clock),
    .reset(Counter_27_reset),
    .io_max(Counter_27_io_max),
    .io_out(Counter_27_io_out),
    .io_enable(Counter_27_io_enable),
    .io_done(Counter_27_io_done)
  );
  Counter_8 Counter_28 (
    .clock(Counter_28_clock),
    .reset(Counter_28_reset),
    .io_max(Counter_28_io_max),
    .io_out(Counter_28_io_out),
    .io_enable(Counter_28_io_enable),
    .io_done(Counter_28_io_done)
  );
  FF_25 FF_74 (
    .clock(FF_74_clock),
    .reset(FF_74_reset),
    .io_in(FF_74_io_in),
    .io_init(FF_74_io_init),
    .io_out(FF_74_io_out),
    .io_enable(FF_74_io_enable)
  );
  Counter_8 Counter_29 (
    .clock(Counter_29_clock),
    .reset(Counter_29_reset),
    .io_max(Counter_29_io_max),
    .io_out(Counter_29_io_out),
    .io_enable(Counter_29_io_enable),
    .io_done(Counter_29_io_done)
  );
  Counter_8 Counter_30 (
    .clock(Counter_30_clock),
    .reset(Counter_30_reset),
    .io_max(Counter_30_io_max),
    .io_out(Counter_30_io_out),
    .io_enable(Counter_30_io_enable),
    .io_done(Counter_30_io_done)
  );
  Counter_8 Counter_31 (
    .clock(Counter_31_clock),
    .reset(Counter_31_reset),
    .io_max(Counter_31_io_max),
    .io_out(Counter_31_io_out),
    .io_enable(Counter_31_io_enable),
    .io_done(Counter_31_io_done)
  );
  Counter_8 Counter_32 (
    .clock(Counter_32_clock),
    .reset(Counter_32_reset),
    .io_max(Counter_32_io_max),
    .io_out(Counter_32_io_out),
    .io_enable(Counter_32_io_enable),
    .io_done(Counter_32_io_done)
  );
  Counter_8 Counter_33 (
    .clock(Counter_33_clock),
    .reset(Counter_33_reset),
    .io_max(Counter_33_io_max),
    .io_out(Counter_33_io_out),
    .io_enable(Counter_33_io_enable),
    .io_done(Counter_33_io_done)
  );
  Counter_8 Counter_34 (
    .clock(Counter_34_clock),
    .reset(Counter_34_reset),
    .io_max(Counter_34_io_max),
    .io_out(Counter_34_io_out),
    .io_enable(Counter_34_io_enable),
    .io_done(Counter_34_io_done)
  );
  Counter_8 Counter_35 (
    .clock(Counter_35_clock),
    .reset(Counter_35_reset),
    .io_max(Counter_35_io_max),
    .io_out(Counter_35_io_out),
    .io_enable(Counter_35_io_enable),
    .io_done(Counter_35_io_done)
  );
  Counter_8 Counter_36 (
    .clock(Counter_36_clock),
    .reset(Counter_36_reset),
    .io_max(Counter_36_io_max),
    .io_out(Counter_36_io_out),
    .io_enable(Counter_36_io_enable),
    .io_done(Counter_36_io_done)
  );
  assign _T_918 = ~ cmdArbiter_io_empty;
  assign _T_919 = io_enable & _T_918;
  assign _T_920 = ~ cmdArbiter_io_deq_0_isWr;
  assign cmdRead = _T_919 & _T_920;
  assign cmdWrite = _T_919 & cmdArbiter_io_deq_0_isWr;
  assign _T_935 = io_dram_cmd_bits_size - 32'h1;
  assign _T_936 = $unsigned(_T_935);
  assign _T_937 = _T_936[31:0];
  assign _T_938 = burstCounter_io_out == _T_937;
  assign _T_939 = wdataMux_io_ins_0_valid & _T_938;
  assign _T_942 = cmdAddr_bits[63:6];
  assign _T_944 = {_T_942,6'h0};
  assign _T_949 = _T_948_bits[15:6];
  assign _T_950 = _T_948_bits[5:0];
  assign _T_952 = _T_950 != 6'h0;
  assign _GEN_0 = {{9'd0}, _T_952};
  assign _T_953 = _T_949 + _GEN_0;
  assign _T_954 = _T_953[9:0];
  assign _T_955 = ~ dramCmdMux_io_out_bits_isWr;
  assign _T_956 = dramCmdMux_io_out_valid & _T_955;
  assign _T_977 = _T_976_bits[15:6];
  assign _T_978 = _T_976_bits[5:0];
  assign _T_980 = _T_978 != 6'h0;
  assign _GEN_1 = {{9'd0}, _T_980};
  assign _T_981 = _T_977 + _GEN_1;
  assign _T_982 = _T_981[9:0];
  assign _T_1035 = io_dram_rresp_bits_tag_streamId == 6'h0;
  assign _T_1036 = io_dram_rresp_valid & _T_1035;
  assign _T_1037 = ~ denseLoadBuffers_0_io_full;
  assign _T_1044 = denseLoadBuffers_0_io_empty & denseLoadBuffers_0_io_deqVld;
  assign _T_1054 = ~ SRFF_sp_io_output_data;
  assign _T_1055 = ~ denseLoadBuffers_0_io_deqVld;
  assign _T_1064 = denseLoadBuffers_0_io_deqVld & _T_1058;
  assign _T_1065 = _T_1054 & _T_1064;
  assign _T_1066 = {denseLoadBuffers_0_io_deq_15,denseLoadBuffers_0_io_deq_14};
  assign _T_1067 = {_T_1066,denseLoadBuffers_0_io_deq_13};
  assign _T_1068 = {_T_1067,denseLoadBuffers_0_io_deq_12};
  assign _T_1069 = {_T_1068,denseLoadBuffers_0_io_deq_11};
  assign _T_1070 = {_T_1069,denseLoadBuffers_0_io_deq_10};
  assign _T_1071 = {_T_1070,denseLoadBuffers_0_io_deq_9};
  assign _T_1072 = {_T_1071,denseLoadBuffers_0_io_deq_8};
  assign _T_1073 = {_T_1072,denseLoadBuffers_0_io_deq_7};
  assign _T_1074 = {_T_1073,denseLoadBuffers_0_io_deq_6};
  assign _T_1075 = {_T_1074,denseLoadBuffers_0_io_deq_5};
  assign _T_1076 = {_T_1075,denseLoadBuffers_0_io_deq_4};
  assign _T_1077 = {_T_1076,denseLoadBuffers_0_io_deq_3};
  assign _T_1078 = {_T_1077,denseLoadBuffers_0_io_deq_2};
  assign _T_1079 = {_T_1078,denseLoadBuffers_0_io_deq_1};
  assign _T_1080 = {_T_1079,denseLoadBuffers_0_io_deq_0};
  assign _T_1084 = ~ SRFF_sp_1_io_output_data;
  assign _T_1085 = ~ denseLoadBuffers_0_io_enqVld;
  assign _T_1094 = denseLoadBuffers_0_io_enqVld & _T_1088;
  assign _T_1095 = _T_1084 & _T_1094;
  assign _T_1096 = {denseLoadBuffers_0_io_enq_15,denseLoadBuffers_0_io_enq_14};
  assign _T_1097 = {_T_1096,denseLoadBuffers_0_io_enq_13};
  assign _T_1098 = {_T_1097,denseLoadBuffers_0_io_enq_12};
  assign _T_1099 = {_T_1098,denseLoadBuffers_0_io_enq_11};
  assign _T_1100 = {_T_1099,denseLoadBuffers_0_io_enq_10};
  assign _T_1101 = {_T_1100,denseLoadBuffers_0_io_enq_9};
  assign _T_1102 = {_T_1101,denseLoadBuffers_0_io_enq_8};
  assign _T_1103 = {_T_1102,denseLoadBuffers_0_io_enq_7};
  assign _T_1104 = {_T_1103,denseLoadBuffers_0_io_enq_6};
  assign _T_1105 = {_T_1104,denseLoadBuffers_0_io_enq_5};
  assign _T_1106 = {_T_1105,denseLoadBuffers_0_io_enq_4};
  assign _T_1107 = {_T_1106,denseLoadBuffers_0_io_enq_3};
  assign _T_1108 = {_T_1107,denseLoadBuffers_0_io_enq_2};
  assign _T_1109 = {_T_1108,denseLoadBuffers_0_io_enq_1};
  assign _T_1110 = {_T_1109,denseLoadBuffers_0_io_enq_0};
  assign _T_1114 = cmdWrite & wdataMux_io_out_valid;
  assign _T_1115 = ~ dramReadySeen;
  assign _T_1116 = _T_1114 & _T_1115;
  assign _T_1117 = ~ denseStoreBuffers_0_io_empty;
  assign _T_1118 = cmdWrite & _T_1117;
  assign _T_1119 = _T_1118 & io_dram_wdata_ready;
  assign _T_1121 = cmdArbiter_io_tag;
  assign _T_1122 = _T_1119 & _T_1121;
  assign _T_1127 = io_dram_wresp_bits_tag_streamId == 6'h1;
  assign _T_1128 = io_dram_wresp_valid & _T_1127;
  assign _T_1129 = ~ FIFOCounter_io_full;
  assign _T_1137 = io_dram_cmd_bits_isWr ? io_dram_cmd_bits_size : 32'h1;
  assign _T_1140 = wdataMux_io_out_valid & io_dram_wdata_ready;
  assign _T_1141 = io_dram_cmd_valid & io_dram_cmd_ready;
  assign _T_1142 = io_dram_cmd_bits_isWr ? _T_1140 : _T_1141;
  assign _T_1150 = io_dram_cmd_valid & io_dram_cmd_bits_isWr;
  assign _T_1151 = burstCounter_io_done | _T_1150;
  assign _T_1153 = io_dram_cmd_ready | dramReadySeen;
  assign _T_1154 = burstCounter_io_done ? 1'h0 : _T_1153;
  assign _T_1160 = io_dram_rresp_valid & io_dram_rresp_ready;
  assign _T_1166 = io_dram_wdata_valid & io_dram_wdata_ready;
  assign _T_1167 = _T_1166 & io_enable;
  assign _T_1173 = io_dram_rresp_ready & io_dram_rresp_valid;
  assign _T_1175 = rdataEnqCount_io_out == 32'h0;
  assign _T_1176 = _T_1173 & _T_1175;
  assign _T_1287 = rdataEnqCount_io_out == 32'h1;
  assign _T_1288 = _T_1173 & _T_1287;
  assign _T_1397 = io_dram_wdata_ready & io_dram_wdata_valid;
  assign _T_1399 = wdataCount_io_out == 32'h0;
  assign _T_1400 = _T_1397 & _T_1399;
  assign _T_1513 = {wdataMux_io_out_bits_wdata_15,wdataMux_io_out_bits_wdata_14};
  assign _T_1514 = {_T_1513,wdataMux_io_out_bits_wdata_13};
  assign _T_1515 = {_T_1514,wdataMux_io_out_bits_wdata_12};
  assign _T_1516 = {_T_1515,wdataMux_io_out_bits_wdata_11};
  assign _T_1517 = {_T_1516,wdataMux_io_out_bits_wdata_10};
  assign _T_1518 = {_T_1517,wdataMux_io_out_bits_wdata_9};
  assign _T_1519 = {_T_1518,wdataMux_io_out_bits_wdata_8};
  assign _T_1520 = {_T_1519,wdataMux_io_out_bits_wdata_7};
  assign _T_1521 = {_T_1520,wdataMux_io_out_bits_wdata_6};
  assign _T_1522 = {_T_1521,wdataMux_io_out_bits_wdata_5};
  assign _T_1523 = {_T_1522,wdataMux_io_out_bits_wdata_4};
  assign _T_1524 = {_T_1523,wdataMux_io_out_bits_wdata_3};
  assign _T_1525 = {_T_1524,wdataMux_io_out_bits_wdata_2};
  assign _T_1526 = {_T_1525,wdataMux_io_out_bits_wdata_1};
  assign _T_1527 = {_T_1526,wdataMux_io_out_bits_wdata_0};
  assign _T_1533 = wdataCount_io_out == 32'h1;
  assign _T_1534 = _T_1397 & _T_1533;
  assign _T_1665 = io_enable & io_dram_cmd_ready;
  assign _T_1666 = _T_1665 & io_dram_cmd_valid;
  assign _T_1674 = io_dram_cmd_ready & io_dram_cmd_valid;
  assign _T_1675 = ~ _T_1674;
  assign _T_1676 = _T_919 & _T_1675;
  assign _T_1685 = _T_1666 & _T_920;
  assign _T_1706 = cmdArbiter_io_tag == 1'h0;
  assign _T_1707 = _T_1141 & _T_1706;
  assign _T_1715 = _T_1666 & cmdArbiter_io_deq_0_isWr;
  assign _T_1737 = _T_1141 & _T_1121;
  assign _T_1749 = io_enable & io_dram_rresp_valid;
  assign _T_1750 = ~ io_dram_rresp_ready;
  assign _T_1751 = _T_1749 & _T_1750;
  assign _T_1757 = ~ io_dram_rresp_valid;
  assign _T_1758 = io_enable & _T_1757;
  assign _T_1759 = _T_1758 & io_dram_rresp_ready;
  assign _T_1768 = _T_1160 & _T_1035;
  assign _T_1774 = io_dram_wresp_valid & io_dram_wresp_ready;
  assign _T_1780 = io_enable & io_dram_wresp_valid;
  assign _T_1781 = ~ io_dram_wresp_ready;
  assign _T_1782 = _T_1780 & _T_1781;
  assign _T_1788 = ~ io_dram_wresp_valid;
  assign _T_1789 = io_enable & _T_1788;
  assign _T_1790 = _T_1789 & io_dram_wresp_ready;
  assign _T_1799 = _T_1774 & _T_1127;
  assign _T_1843 = io_dram_rresp_bits_tag_streamId >= 6'h1;
  assign _T_1872 = io_dram_rresp_valid & denseLoadBuffers_0_io_enqVld;
  assign _T_1885 = _T_1160 & denseLoadBuffers_0_io_enqVld;
  assign _T_1892 = io_dram_rresp_valid & _T_1750;
  assign io_dram_cmd_valid = dramCmdMux_io_out_valid;
  assign io_dram_cmd_bits_addr = dramCmdMux_io_out_bits_addr;
  assign io_dram_cmd_bits_size = dramCmdMux_io_out_bits_size;
  assign io_dram_cmd_bits_isWr = dramCmdMux_io_out_bits_isWr;
  assign io_dram_cmd_bits_tag_uid = dramCmdMux_io_out_bits_tag_uid;
  assign io_dram_cmd_bits_tag_streamId = dramCmdMux_io_out_bits_tag_streamId;
  assign io_dram_wdata_valid = wdataMux_io_out_valid;
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0;
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1;
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2;
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3;
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4;
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5;
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6;
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7;
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8;
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9;
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10;
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11;
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12;
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13;
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14;
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15;
  assign io_dram_wdata_bits_wlast = wdataMux_io_out_bits_wlast;
  assign io_dram_rresp_ready = rrespReadyMux_io_out;
  assign io_dram_wresp_ready = wrespReadyMux_io_out;
  assign io_debugSignals_0 = {{26'd0}, FF_io_out};
  assign io_debugSignals_1 = FF_1_io_out[31:0];
  assign io_debugSignals_2 = FF_2_io_out;
  assign io_debugSignals_3 = {{31'd0}, FF_3_io_out};
  assign io_debugSignals_4 = FF_4_io_out[31:0];
  assign io_debugSignals_5 = {{16'd0}, FF_5_io_out};
  assign io_debugSignals_6 = Counter_io_out;
  assign io_debugSignals_7 = Counter_1_io_out;
  assign io_debugSignals_8 = FF_6_io_out[31:0];
  assign io_debugSignals_9 = FF_7_io_out[31:0];
  assign io_debugSignals_10 = Counter_2_io_out;
  assign io_debugSignals_11 = cycleCount_io_out;
  assign io_debugSignals_12 = FF_8_io_out;
  assign io_debugSignals_13 = FF_9_io_out;
  assign io_debugSignals_14 = FF_10_io_out;
  assign io_debugSignals_15 = FF_11_io_out;
  assign io_debugSignals_16 = FF_12_io_out;
  assign io_debugSignals_17 = FF_13_io_out;
  assign io_debugSignals_18 = FF_14_io_out;
  assign io_debugSignals_19 = FF_15_io_out;
  assign io_debugSignals_20 = FF_16_io_out;
  assign io_debugSignals_21 = FF_17_io_out;
  assign io_debugSignals_22 = FF_18_io_out;
  assign io_debugSignals_23 = FF_19_io_out;
  assign io_debugSignals_24 = FF_20_io_out;
  assign io_debugSignals_25 = FF_21_io_out;
  assign io_debugSignals_26 = FF_22_io_out;
  assign io_debugSignals_27 = FF_23_io_out;
  assign io_debugSignals_28 = FF_24_io_out;
  assign io_debugSignals_29 = FF_25_io_out;
  assign io_debugSignals_30 = FF_26_io_out;
  assign io_debugSignals_31 = FF_27_io_out;
  assign io_debugSignals_32 = FF_28_io_out;
  assign io_debugSignals_33 = FF_29_io_out;
  assign io_debugSignals_34 = FF_30_io_out;
  assign io_debugSignals_35 = FF_31_io_out;
  assign io_debugSignals_36 = FF_32_io_out;
  assign io_debugSignals_37 = FF_33_io_out;
  assign io_debugSignals_38 = FF_34_io_out;
  assign io_debugSignals_39 = FF_35_io_out;
  assign io_debugSignals_40 = FF_36_io_out;
  assign io_debugSignals_41 = FF_37_io_out;
  assign io_debugSignals_42 = FF_38_io_out;
  assign io_debugSignals_43 = FF_39_io_out;
  assign io_debugSignals_44 = FF_40_io_out;
  assign io_debugSignals_45 = FF_41_io_out;
  assign io_debugSignals_46 = FF_42_io_out;
  assign io_debugSignals_47 = FF_43_io_out;
  assign io_debugSignals_48 = FF_44_io_out;
  assign io_debugSignals_49 = FF_45_io_out;
  assign io_debugSignals_50 = FF_46_io_out;
  assign io_debugSignals_51 = FF_47_io_out;
  assign io_debugSignals_52 = FF_48_io_out;
  assign io_debugSignals_53 = FF_49_io_out;
  assign io_debugSignals_54 = FF_50_io_out;
  assign io_debugSignals_55 = FF_51_io_out;
  assign io_debugSignals_56 = FF_52_io_out;
  assign io_debugSignals_57 = FF_53_io_out;
  assign io_debugSignals_58 = FF_54_io_out;
  assign io_debugSignals_59 = FF_55_io_out;
  assign io_debugSignals_60 = FF_56_io_out[31:0];
  assign io_debugSignals_61 = FF_57_io_out;
  assign io_debugSignals_62 = FF_58_io_out;
  assign io_debugSignals_63 = FF_59_io_out;
  assign io_debugSignals_64 = FF_60_io_out;
  assign io_debugSignals_65 = FF_61_io_out;
  assign io_debugSignals_66 = FF_62_io_out;
  assign io_debugSignals_67 = FF_63_io_out;
  assign io_debugSignals_68 = FF_64_io_out;
  assign io_debugSignals_69 = FF_65_io_out;
  assign io_debugSignals_70 = FF_66_io_out;
  assign io_debugSignals_71 = FF_67_io_out;
  assign io_debugSignals_72 = FF_68_io_out;
  assign io_debugSignals_73 = FF_69_io_out;
  assign io_debugSignals_74 = FF_70_io_out;
  assign io_debugSignals_75 = FF_71_io_out;
  assign io_debugSignals_76 = FF_72_io_out;
  assign io_debugSignals_77 = FF_73_io_out[31:0];
  assign io_debugSignals_78 = Counter_3_io_out;
  assign io_debugSignals_79 = Counter_4_io_out;
  assign io_debugSignals_80 = Counter_5_io_out;
  assign io_debugSignals_81 = Counter_7_io_out;
  assign io_debugSignals_82 = Counter_8_io_out;
  assign io_debugSignals_83 = Counter_6_io_out;
  assign io_debugSignals_84 = Counter_9_io_out;
  assign io_debugSignals_85 = Counter_11_io_out;
  assign io_debugSignals_86 = Counter_12_io_out;
  assign io_debugSignals_87 = Counter_10_io_out;
  assign io_debugSignals_88 = Counter_13_io_out;
  assign io_debugSignals_89 = Counter_14_io_out;
  assign io_debugSignals_90 = Counter_15_io_out;
  assign io_debugSignals_91 = Counter_16_io_out;
  assign io_debugSignals_92 = Counter_17_io_out;
  assign io_debugSignals_93 = Counter_18_io_out;
  assign io_debugSignals_94 = Counter_19_io_out;
  assign io_debugSignals_95 = Counter_20_io_out;
  assign io_debugSignals_96 = Counter_21_io_out;
  assign io_debugSignals_97 = Counter_22_io_out;
  assign io_debugSignals_98 = Counter_23_io_out;
  assign io_debugSignals_99 = Counter_24_io_out;
  assign io_debugSignals_100 = Counter_25_io_out;
  assign io_debugSignals_101 = Counter_26_io_out;
  assign io_debugSignals_102 = Counter_27_io_out;
  assign io_debugSignals_103 = Counter_28_io_out;
  assign io_debugSignals_104 = {{26'd0}, FF_74_io_out};
  assign io_debugSignals_105 = Counter_29_io_out;
  assign io_debugSignals_106 = Counter_30_io_out;
  assign io_debugSignals_107 = Counter_31_io_out;
  assign io_debugSignals_108 = Counter_32_io_out;
  assign io_debugSignals_109 = Counter_33_io_out;
  assign io_debugSignals_110 = Counter_34_io_out;
  assign io_debugSignals_111 = Counter_35_io_out;
  assign io_debugSignals_112 = Counter_36_io_out;
  assign io_debugSignals_113 = wdataCount_io_out;
  assign cmdArbiter_io_fifo_0_deq_0_addr = cmdFifos_0_io_deq_0_addr;
  assign cmdArbiter_io_fifo_0_deq_0_isWr = cmdFifos_0_io_deq_0_isWr;
  assign cmdArbiter_io_fifo_0_deq_0_size = cmdFifos_0_io_deq_0_size;
  assign cmdArbiter_io_fifo_0_empty = cmdFifos_0_io_empty;
  assign cmdArbiter_io_fifo_0_almostEmpty = cmdFifos_0_io_almostEmpty;
  assign cmdArbiter_io_fifo_1_deq_0_addr = cmdFifos_1_io_deq_0_addr;
  assign cmdArbiter_io_fifo_1_deq_0_isWr = cmdFifos_1_io_deq_0_isWr;
  assign cmdArbiter_io_fifo_1_deq_0_size = cmdFifos_1_io_deq_0_size;
  assign cmdArbiter_io_fifo_1_empty = cmdFifos_1_io_empty;
  assign cmdArbiter_io_deqVld = cmdDeqValidMux_io_out;
  assign cmdArbiter_clock = clock;
  assign cmdArbiter_reset = reset;
  assign cmdFifos_0_io_deqVld = cmdArbiter_io_fifo_0_deqVld;
  assign cmdFifos_0_clock = clock;
  assign cmdFifos_0_reset = reset;
  assign cmdFifos_1_io_deqVld = cmdArbiter_io_fifo_1_deqVld;
  assign cmdFifos_1_clock = clock;
  assign cmdFifos_1_reset = reset;
  assign cmdAddr_bits = cmdArbiter_io_deq_0_addr;
  assign burstCounter_io_max = _T_1137;
  assign burstCounter_io_enable = _T_1142;
  assign burstCounter_clock = clock;
  assign burstCounter_reset = reset;
  assign burstTagCounter_io_max = 10'h3ff;
  assign burstTagCounter_io_enable = _T_1141;
  assign burstTagCounter_clock = clock;
  assign burstTagCounter_reset = reset;
  assign dramReadySeen = dramReadyFF_io_out;
  assign rrespReadyMux_io_ins_0 = _T_1037;
  assign wdataMux_io_ins_0_valid = _T_1118;
  assign wdataMux_io_ins_0_bits_wdata_0 = denseStoreBuffers_0_io_deq_0;
  assign wdataMux_io_ins_0_bits_wdata_1 = denseStoreBuffers_0_io_deq_1;
  assign wdataMux_io_ins_0_bits_wdata_2 = denseStoreBuffers_0_io_deq_2;
  assign wdataMux_io_ins_0_bits_wdata_3 = denseStoreBuffers_0_io_deq_3;
  assign wdataMux_io_ins_0_bits_wdata_4 = denseStoreBuffers_0_io_deq_4;
  assign wdataMux_io_ins_0_bits_wdata_5 = denseStoreBuffers_0_io_deq_5;
  assign wdataMux_io_ins_0_bits_wdata_6 = denseStoreBuffers_0_io_deq_6;
  assign wdataMux_io_ins_0_bits_wdata_7 = denseStoreBuffers_0_io_deq_7;
  assign wdataMux_io_ins_0_bits_wdata_8 = denseStoreBuffers_0_io_deq_8;
  assign wdataMux_io_ins_0_bits_wdata_9 = denseStoreBuffers_0_io_deq_9;
  assign wdataMux_io_ins_0_bits_wdata_10 = denseStoreBuffers_0_io_deq_10;
  assign wdataMux_io_ins_0_bits_wdata_11 = denseStoreBuffers_0_io_deq_11;
  assign wdataMux_io_ins_0_bits_wdata_12 = denseStoreBuffers_0_io_deq_12;
  assign wdataMux_io_ins_0_bits_wdata_13 = denseStoreBuffers_0_io_deq_13;
  assign wdataMux_io_ins_0_bits_wdata_14 = denseStoreBuffers_0_io_deq_14;
  assign wdataMux_io_ins_0_bits_wdata_15 = denseStoreBuffers_0_io_deq_15;
  assign wdataMux_io_ins_0_bits_wlast = _T_939;
  assign cmdDeqValidMux_io_ins_0 = io_dram_cmd_ready;
  assign cmdDeqValidMux_io_ins_1 = burstCounter_io_done;
  assign cmdDeqValidMux_io_sel = cmdArbiter_io_tag;
  assign dramCmdMux_io_ins_0_valid = cmdRead;
  assign dramCmdMux_io_ins_0_bits_addr = _T_944;
  assign dramCmdMux_io_ins_0_bits_size = {{22'd0}, _T_954};
  assign dramCmdMux_io_ins_0_bits_isWr = cmdArbiter_io_deq_0_isWr;
  assign dramCmdMux_io_ins_0_bits_tag_uid = {{16'd0}, burstTagCounter_io_out};
  assign dramCmdMux_io_ins_0_bits_tag_streamId = _T_946_streamId;
  assign dramCmdMux_io_ins_1_valid = _T_1116;
  assign dramCmdMux_io_ins_1_bits_addr = _T_944;
  assign dramCmdMux_io_ins_1_bits_size = {{22'd0}, _T_982};
  assign dramCmdMux_io_ins_1_bits_isWr = cmdArbiter_io_deq_0_isWr;
  assign dramCmdMux_io_ins_1_bits_tag_uid = {{16'd0}, burstTagCounter_io_out};
  assign dramCmdMux_io_ins_1_bits_tag_streamId = _T_974_streamId;
  assign dramCmdMux_io_sel = cmdArbiter_io_tag;
  assign _T_946_streamId = {{5'd0}, cmdArbiter_io_tag};
  assign _T_948_bits = cmdArbiter_io_deq_0_size;
  assign FF_io_in = dramCmdMux_io_out_bits_tag_streamId;
  assign FF_io_init = 6'h3e;
  assign FF_io_enable = _T_956;
  assign FF_clock = clock;
  assign FF_reset = reset;
  assign FF_1_io_in = dramCmdMux_io_out_bits_addr;
  assign FF_1_io_init = 64'h175bf;
  assign FF_1_io_enable = _T_956;
  assign FF_1_clock = clock;
  assign FF_1_reset = reset;
  assign FF_2_io_in = dramCmdMux_io_out_bits_size;
  assign FF_2_io_init = 32'h2eb7e;
  assign FF_2_io_enable = _T_956;
  assign FF_2_clock = clock;
  assign FF_2_reset = reset;
  assign _T_974_streamId = {{5'd0}, cmdArbiter_io_tag};
  assign _T_976_bits = cmdArbiter_io_deq_0_size;
  assign FF_3_io_in = cmdArbiter_io_tag;
  assign FF_3_io_init = 1'h1;
  assign FF_3_io_enable = cmdWrite;
  assign FF_3_clock = clock;
  assign FF_3_reset = reset;
  assign FF_4_io_in = cmdAddr_bits;
  assign FF_4_io_init = 64'h5d6fc;
  assign FF_4_io_enable = cmdWrite;
  assign FF_4_clock = clock;
  assign FF_4_reset = reset;
  assign FF_5_io_in = cmdArbiter_io_deq_0_size;
  assign FF_5_io_enable = cmdWrite;
  assign FF_5_clock = clock;
  assign FF_5_reset = reset;
  assign wrespReadyMux_io_ins_0 = _T_1129;
  assign gatherLoadIssueMux_io_ins_0 = 1'h0;
  assign gatherLoadIssueMux_io_ins_1 = 1'h0;
  assign gatherLoadIssueMux_io_sel = cmdArbiter_io_tag;
  assign gatherLoadIssue_io_max = 32'hffffffff;
  assign gatherLoadIssue_io_enable = gatherLoadIssueMux_io_out;
  assign gatherLoadIssue_clock = clock;
  assign gatherLoadIssue_reset = reset;
  assign gatherLoadSkipMux_io_ins_0 = 1'h0;
  assign gatherLoadSkipMux_io_ins_1 = 1'h0;
  assign gatherLoadSkipMux_io_sel = cmdArbiter_io_tag;
  assign gatherLoadSkip_io_max = 32'hffffffff;
  assign gatherLoadSkip_io_enable = gatherLoadSkipMux_io_out;
  assign gatherLoadSkip_clock = clock;
  assign gatherLoadSkip_reset = reset;
  assign scatterLoadIssueMux_io_ins_0 = 1'h0;
  assign scatterLoadIssueMux_io_ins_1 = 1'h0;
  assign scatterLoadIssueMux_io_sel = cmdArbiter_io_tag;
  assign scatterLoadIssue_io_max = 32'hffffffff;
  assign scatterLoadIssue_io_enable = scatterLoadIssueMux_io_out;
  assign scatterLoadIssue_clock = clock;
  assign scatterLoadIssue_reset = reset;
  assign scatterLoadSkipMux_io_ins_0 = 1'h0;
  assign scatterLoadSkipMux_io_ins_1 = 1'h0;
  assign scatterLoadSkipMux_io_sel = cmdArbiter_io_tag;
  assign scatterLoadSkip_io_max = 32'hffffffff;
  assign scatterLoadSkip_io_enable = scatterLoadSkipMux_io_out;
  assign scatterLoadSkip_clock = clock;
  assign scatterLoadSkip_reset = reset;
  assign scatterStoreIssueMux_io_ins_0 = 1'h0;
  assign scatterStoreIssueMux_io_ins_1 = 1'h0;
  assign scatterStoreIssueMux_io_sel = cmdArbiter_io_tag;
  assign scatterStoreIssue_io_max = 32'hffffffff;
  assign scatterStoreIssue_io_enable = scatterStoreIssueMux_io_out;
  assign scatterStoreIssue_clock = clock;
  assign scatterStoreIssue_reset = reset;
  assign scatterStoreSkipMux_io_ins_0 = 1'h0;
  assign scatterStoreSkipMux_io_ins_1 = 1'h0;
  assign scatterStoreSkipMux_io_sel = cmdArbiter_io_tag;
  assign scatterStoreSkip_io_max = 32'hffffffff;
  assign scatterStoreSkip_io_enable = scatterStoreSkipMux_io_out;
  assign scatterStoreSkip_clock = clock;
  assign scatterStoreSkip_reset = reset;
  assign denseLoadBuffers_0_io_enq_0 = io_dram_rresp_bits_rdata_0;
  assign denseLoadBuffers_0_io_enq_1 = io_dram_rresp_bits_rdata_1;
  assign denseLoadBuffers_0_io_enq_2 = io_dram_rresp_bits_rdata_2;
  assign denseLoadBuffers_0_io_enq_3 = io_dram_rresp_bits_rdata_3;
  assign denseLoadBuffers_0_io_enq_4 = io_dram_rresp_bits_rdata_4;
  assign denseLoadBuffers_0_io_enq_5 = io_dram_rresp_bits_rdata_5;
  assign denseLoadBuffers_0_io_enq_6 = io_dram_rresp_bits_rdata_6;
  assign denseLoadBuffers_0_io_enq_7 = io_dram_rresp_bits_rdata_7;
  assign denseLoadBuffers_0_io_enq_8 = io_dram_rresp_bits_rdata_8;
  assign denseLoadBuffers_0_io_enq_9 = io_dram_rresp_bits_rdata_9;
  assign denseLoadBuffers_0_io_enq_10 = io_dram_rresp_bits_rdata_10;
  assign denseLoadBuffers_0_io_enq_11 = io_dram_rresp_bits_rdata_11;
  assign denseLoadBuffers_0_io_enq_12 = io_dram_rresp_bits_rdata_12;
  assign denseLoadBuffers_0_io_enq_13 = io_dram_rresp_bits_rdata_13;
  assign denseLoadBuffers_0_io_enq_14 = io_dram_rresp_bits_rdata_14;
  assign denseLoadBuffers_0_io_enq_15 = io_dram_rresp_bits_rdata_15;
  assign denseLoadBuffers_0_io_enqVld = _T_1036;
  assign denseLoadBuffers_0_io_deqVld = 1'h0;
  assign denseLoadBuffers_0_clock = clock;
  assign denseLoadBuffers_0_reset = reset;
  assign Counter_io_max = 32'hffffffff;
  assign Counter_io_enable = denseLoadBuffers_0_io_enqVld;
  assign Counter_clock = clock;
  assign Counter_reset = reset;
  assign Counter_1_io_max = 32'hffffffff;
  assign Counter_1_io_enable = _T_1044;
  assign Counter_1_clock = clock;
  assign Counter_1_reset = reset;
  assign SRFF_sp_io_input_set = denseLoadBuffers_0_io_deqVld;
  assign SRFF_sp_io_input_reset = reset;
  assign SRFF_sp_io_input_asyn_reset = reset;
  assign SRFF_sp_clock = clock;
  assign SRFF_sp_reset = reset;
  assign SRFF_sp_1_io_input_set = denseLoadBuffers_0_io_enqVld;
  assign SRFF_sp_1_io_input_reset = reset;
  assign SRFF_sp_1_io_input_asyn_reset = reset;
  assign SRFF_sp_1_clock = clock;
  assign SRFF_sp_1_reset = reset;
  assign FF_6_io_in = _T_1080;
  assign FF_6_io_init = 512'hbadf8;
  assign FF_6_io_enable = _T_1065;
  assign FF_6_clock = clock;
  assign FF_6_reset = reset;
  assign FF_7_io_in = _T_1110;
  assign FF_7_io_init = 512'hbadf9;
  assign FF_7_io_enable = _T_1095;
  assign FF_7_clock = clock;
  assign FF_7_reset = reset;
  assign denseStoreBuffers_0_io_enq_0 = 32'h0;
  assign denseStoreBuffers_0_io_enq_1 = 32'h0;
  assign denseStoreBuffers_0_io_enq_2 = 32'h0;
  assign denseStoreBuffers_0_io_enq_3 = 32'h0;
  assign denseStoreBuffers_0_io_enq_4 = 32'h0;
  assign denseStoreBuffers_0_io_enq_5 = 32'h0;
  assign denseStoreBuffers_0_io_enq_6 = 32'h0;
  assign denseStoreBuffers_0_io_enq_7 = 32'h0;
  assign denseStoreBuffers_0_io_enq_8 = 32'h0;
  assign denseStoreBuffers_0_io_enq_9 = 32'h0;
  assign denseStoreBuffers_0_io_enq_10 = 32'h0;
  assign denseStoreBuffers_0_io_enq_11 = 32'h0;
  assign denseStoreBuffers_0_io_enq_12 = 32'h0;
  assign denseStoreBuffers_0_io_enq_13 = 32'h0;
  assign denseStoreBuffers_0_io_enq_14 = 32'h0;
  assign denseStoreBuffers_0_io_enq_15 = 32'h0;
  assign denseStoreBuffers_0_io_enqVld = 1'h0;
  assign denseStoreBuffers_0_io_deqVld = _T_1122;
  assign denseStoreBuffers_0_clock = clock;
  assign denseStoreBuffers_0_reset = reset;
  assign FIFOCounter_io_enqVld = _T_1128;
  assign FIFOCounter_clock = clock;
  assign FIFOCounter_reset = reset;
  assign Counter_2_io_max = 32'hffffffff;
  assign Counter_2_io_enable = FIFOCounter_io_enqVld;
  assign Counter_2_clock = clock;
  assign Counter_2_reset = reset;
  assign dramReadyFF_io_in = _T_1154;
  assign dramReadyFF_io_init = 1'h0;
  assign dramReadyFF_io_enable = _T_1151;
  assign dramReadyFF_clock = clock;
  assign dramReadyFF_reset = reset;
  assign cycleCount_io_max = 32'hffffffff;
  assign cycleCount_io_enable = io_enable;
  assign cycleCount_clock = clock;
  assign cycleCount_reset = reset;
  assign rdataEnqCount_io_max = 32'hffffffff;
  assign rdataEnqCount_io_enable = _T_1160;
  assign rdataEnqCount_clock = clock;
  assign rdataEnqCount_reset = reset;
  assign wdataCount_io_max = 32'hffffffff;
  assign wdataCount_io_enable = _T_1167;
  assign wdataCount_clock = clock;
  assign wdataCount_reset = reset;
  assign FF_8_io_in = io_dram_rresp_bits_rdata_0;
  assign FF_8_io_init = 32'hbadfc;
  assign FF_8_io_enable = _T_1176;
  assign FF_8_clock = clock;
  assign FF_8_reset = reset;
  assign FF_9_io_in = io_dram_rresp_bits_rdata_1;
  assign FF_9_io_init = 32'hbadfd;
  assign FF_9_io_enable = _T_1176;
  assign FF_9_clock = clock;
  assign FF_9_reset = reset;
  assign FF_10_io_in = io_dram_rresp_bits_rdata_2;
  assign FF_10_io_init = 32'hbadfe;
  assign FF_10_io_enable = _T_1176;
  assign FF_10_clock = clock;
  assign FF_10_reset = reset;
  assign FF_11_io_in = io_dram_rresp_bits_rdata_3;
  assign FF_11_io_init = 32'hbadff;
  assign FF_11_io_enable = _T_1176;
  assign FF_11_clock = clock;
  assign FF_11_reset = reset;
  assign FF_12_io_in = io_dram_rresp_bits_rdata_4;
  assign FF_12_io_init = 32'h175bf0;
  assign FF_12_io_enable = _T_1176;
  assign FF_12_clock = clock;
  assign FF_12_reset = reset;
  assign FF_13_io_in = io_dram_rresp_bits_rdata_5;
  assign FF_13_io_init = 32'h175bf1;
  assign FF_13_io_enable = _T_1176;
  assign FF_13_clock = clock;
  assign FF_13_reset = reset;
  assign FF_14_io_in = io_dram_rresp_bits_rdata_6;
  assign FF_14_io_init = 32'h175bf2;
  assign FF_14_io_enable = _T_1176;
  assign FF_14_clock = clock;
  assign FF_14_reset = reset;
  assign FF_15_io_in = io_dram_rresp_bits_rdata_7;
  assign FF_15_io_init = 32'h175bf3;
  assign FF_15_io_enable = _T_1176;
  assign FF_15_clock = clock;
  assign FF_15_reset = reset;
  assign FF_16_io_in = io_dram_rresp_bits_rdata_8;
  assign FF_16_io_init = 32'h175bf4;
  assign FF_16_io_enable = _T_1176;
  assign FF_16_clock = clock;
  assign FF_16_reset = reset;
  assign FF_17_io_in = io_dram_rresp_bits_rdata_9;
  assign FF_17_io_init = 32'h175bf5;
  assign FF_17_io_enable = _T_1176;
  assign FF_17_clock = clock;
  assign FF_17_reset = reset;
  assign FF_18_io_in = io_dram_rresp_bits_rdata_10;
  assign FF_18_io_init = 32'h175bf6;
  assign FF_18_io_enable = _T_1176;
  assign FF_18_clock = clock;
  assign FF_18_reset = reset;
  assign FF_19_io_in = io_dram_rresp_bits_rdata_11;
  assign FF_19_io_init = 32'h175bf7;
  assign FF_19_io_enable = _T_1176;
  assign FF_19_clock = clock;
  assign FF_19_reset = reset;
  assign FF_20_io_in = io_dram_rresp_bits_rdata_12;
  assign FF_20_io_init = 32'h175bf8;
  assign FF_20_io_enable = _T_1176;
  assign FF_20_clock = clock;
  assign FF_20_reset = reset;
  assign FF_21_io_in = io_dram_rresp_bits_rdata_13;
  assign FF_21_io_init = 32'h175bf9;
  assign FF_21_io_enable = _T_1176;
  assign FF_21_clock = clock;
  assign FF_21_reset = reset;
  assign FF_22_io_in = io_dram_rresp_bits_rdata_14;
  assign FF_22_io_init = 32'h175bfa;
  assign FF_22_io_enable = _T_1176;
  assign FF_22_clock = clock;
  assign FF_22_reset = reset;
  assign FF_23_io_in = io_dram_rresp_bits_rdata_15;
  assign FF_23_io_init = 32'h175bfb;
  assign FF_23_io_enable = _T_1176;
  assign FF_23_clock = clock;
  assign FF_23_reset = reset;
  assign FF_24_io_in = io_dram_rresp_bits_rdata_0;
  assign FF_24_io_init = 32'h175bfc;
  assign FF_24_io_enable = _T_1288;
  assign FF_24_clock = clock;
  assign FF_24_reset = reset;
  assign FF_25_io_in = io_dram_rresp_bits_rdata_1;
  assign FF_25_io_init = 32'h175bfd;
  assign FF_25_io_enable = _T_1288;
  assign FF_25_clock = clock;
  assign FF_25_reset = reset;
  assign FF_26_io_in = io_dram_rresp_bits_rdata_2;
  assign FF_26_io_init = 32'h175bfe;
  assign FF_26_io_enable = _T_1288;
  assign FF_26_clock = clock;
  assign FF_26_reset = reset;
  assign FF_27_io_in = io_dram_rresp_bits_rdata_3;
  assign FF_27_io_init = 32'h175bff;
  assign FF_27_io_enable = _T_1288;
  assign FF_27_clock = clock;
  assign FF_27_reset = reset;
  assign FF_28_io_in = io_dram_rresp_bits_rdata_4;
  assign FF_28_io_init = 32'h2eb7e0;
  assign FF_28_io_enable = _T_1288;
  assign FF_28_clock = clock;
  assign FF_28_reset = reset;
  assign FF_29_io_in = io_dram_rresp_bits_rdata_5;
  assign FF_29_io_init = 32'h2eb7e1;
  assign FF_29_io_enable = _T_1288;
  assign FF_29_clock = clock;
  assign FF_29_reset = reset;
  assign FF_30_io_in = io_dram_rresp_bits_rdata_6;
  assign FF_30_io_init = 32'h2eb7e2;
  assign FF_30_io_enable = _T_1288;
  assign FF_30_clock = clock;
  assign FF_30_reset = reset;
  assign FF_31_io_in = io_dram_rresp_bits_rdata_7;
  assign FF_31_io_init = 32'h2eb7e3;
  assign FF_31_io_enable = _T_1288;
  assign FF_31_clock = clock;
  assign FF_31_reset = reset;
  assign FF_32_io_in = io_dram_rresp_bits_rdata_8;
  assign FF_32_io_init = 32'h2eb7e4;
  assign FF_32_io_enable = _T_1288;
  assign FF_32_clock = clock;
  assign FF_32_reset = reset;
  assign FF_33_io_in = io_dram_rresp_bits_rdata_9;
  assign FF_33_io_init = 32'h2eb7e5;
  assign FF_33_io_enable = _T_1288;
  assign FF_33_clock = clock;
  assign FF_33_reset = reset;
  assign FF_34_io_in = io_dram_rresp_bits_rdata_10;
  assign FF_34_io_init = 32'h2eb7e6;
  assign FF_34_io_enable = _T_1288;
  assign FF_34_clock = clock;
  assign FF_34_reset = reset;
  assign FF_35_io_in = io_dram_rresp_bits_rdata_11;
  assign FF_35_io_init = 32'h2eb7e7;
  assign FF_35_io_enable = _T_1288;
  assign FF_35_clock = clock;
  assign FF_35_reset = reset;
  assign FF_36_io_in = io_dram_rresp_bits_rdata_12;
  assign FF_36_io_init = 32'h2eb7e8;
  assign FF_36_io_enable = _T_1288;
  assign FF_36_clock = clock;
  assign FF_36_reset = reset;
  assign FF_37_io_in = io_dram_rresp_bits_rdata_13;
  assign FF_37_io_init = 32'h2eb7e9;
  assign FF_37_io_enable = _T_1288;
  assign FF_37_clock = clock;
  assign FF_37_reset = reset;
  assign FF_38_io_in = io_dram_rresp_bits_rdata_14;
  assign FF_38_io_init = 32'h2eb7ea;
  assign FF_38_io_enable = _T_1288;
  assign FF_38_clock = clock;
  assign FF_38_reset = reset;
  assign FF_39_io_in = io_dram_rresp_bits_rdata_15;
  assign FF_39_io_init = 32'h2eb7eb;
  assign FF_39_io_enable = _T_1288;
  assign FF_39_clock = clock;
  assign FF_39_reset = reset;
  assign FF_40_io_in = io_dram_wdata_bits_wdata_0;
  assign FF_40_io_init = 32'h2eb7ec;
  assign FF_40_io_enable = _T_1400;
  assign FF_40_clock = clock;
  assign FF_40_reset = reset;
  assign FF_41_io_in = io_dram_wdata_bits_wdata_1;
  assign FF_41_io_init = 32'h2eb7ed;
  assign FF_41_io_enable = _T_1400;
  assign FF_41_clock = clock;
  assign FF_41_reset = reset;
  assign FF_42_io_in = io_dram_wdata_bits_wdata_2;
  assign FF_42_io_init = 32'h2eb7ee;
  assign FF_42_io_enable = _T_1400;
  assign FF_42_clock = clock;
  assign FF_42_reset = reset;
  assign FF_43_io_in = io_dram_wdata_bits_wdata_3;
  assign FF_43_io_init = 32'h2eb7ef;
  assign FF_43_io_enable = _T_1400;
  assign FF_43_clock = clock;
  assign FF_43_reset = reset;
  assign FF_44_io_in = io_dram_wdata_bits_wdata_4;
  assign FF_44_io_init = 32'h2eb7f0;
  assign FF_44_io_enable = _T_1400;
  assign FF_44_clock = clock;
  assign FF_44_reset = reset;
  assign FF_45_io_in = io_dram_wdata_bits_wdata_5;
  assign FF_45_io_init = 32'h2eb7f1;
  assign FF_45_io_enable = _T_1400;
  assign FF_45_clock = clock;
  assign FF_45_reset = reset;
  assign FF_46_io_in = io_dram_wdata_bits_wdata_6;
  assign FF_46_io_init = 32'h2eb7f2;
  assign FF_46_io_enable = _T_1400;
  assign FF_46_clock = clock;
  assign FF_46_reset = reset;
  assign FF_47_io_in = io_dram_wdata_bits_wdata_7;
  assign FF_47_io_init = 32'h2eb7f3;
  assign FF_47_io_enable = _T_1400;
  assign FF_47_clock = clock;
  assign FF_47_reset = reset;
  assign FF_48_io_in = io_dram_wdata_bits_wdata_8;
  assign FF_48_io_init = 32'h2eb7f4;
  assign FF_48_io_enable = _T_1400;
  assign FF_48_clock = clock;
  assign FF_48_reset = reset;
  assign FF_49_io_in = io_dram_wdata_bits_wdata_9;
  assign FF_49_io_init = 32'h2eb7f5;
  assign FF_49_io_enable = _T_1400;
  assign FF_49_clock = clock;
  assign FF_49_reset = reset;
  assign FF_50_io_in = io_dram_wdata_bits_wdata_10;
  assign FF_50_io_init = 32'h2eb7f6;
  assign FF_50_io_enable = _T_1400;
  assign FF_50_clock = clock;
  assign FF_50_reset = reset;
  assign FF_51_io_in = io_dram_wdata_bits_wdata_11;
  assign FF_51_io_init = 32'h2eb7f7;
  assign FF_51_io_enable = _T_1400;
  assign FF_51_clock = clock;
  assign FF_51_reset = reset;
  assign FF_52_io_in = io_dram_wdata_bits_wdata_12;
  assign FF_52_io_init = 32'h2eb7f8;
  assign FF_52_io_enable = _T_1400;
  assign FF_52_clock = clock;
  assign FF_52_reset = reset;
  assign FF_53_io_in = io_dram_wdata_bits_wdata_13;
  assign FF_53_io_init = 32'h2eb7f9;
  assign FF_53_io_enable = _T_1400;
  assign FF_53_clock = clock;
  assign FF_53_reset = reset;
  assign FF_54_io_in = io_dram_wdata_bits_wdata_14;
  assign FF_54_io_init = 32'h2eb7fa;
  assign FF_54_io_enable = _T_1400;
  assign FF_54_clock = clock;
  assign FF_54_reset = reset;
  assign FF_55_io_in = io_dram_wdata_bits_wdata_15;
  assign FF_55_io_init = 32'h2eb7fb;
  assign FF_55_io_enable = _T_1400;
  assign FF_55_clock = clock;
  assign FF_55_reset = reset;
  assign FF_56_io_in = _T_1527;
  assign FF_56_io_init = 512'h2eb7fc;
  assign FF_56_io_enable = _T_1400;
  assign FF_56_clock = clock;
  assign FF_56_reset = reset;
  assign FF_57_io_in = io_dram_wdata_bits_wdata_0;
  assign FF_57_io_init = 32'h2eb7fd;
  assign FF_57_io_enable = _T_1534;
  assign FF_57_clock = clock;
  assign FF_57_reset = reset;
  assign FF_58_io_in = io_dram_wdata_bits_wdata_1;
  assign FF_58_io_init = 32'h2eb7fe;
  assign FF_58_io_enable = _T_1534;
  assign FF_58_clock = clock;
  assign FF_58_reset = reset;
  assign FF_59_io_in = io_dram_wdata_bits_wdata_2;
  assign FF_59_io_init = 32'h2eb7ff;
  assign FF_59_io_enable = _T_1534;
  assign FF_59_clock = clock;
  assign FF_59_reset = reset;
  assign FF_60_io_in = io_dram_wdata_bits_wdata_3;
  assign FF_60_io_init = 32'h5d6fc0;
  assign FF_60_io_enable = _T_1534;
  assign FF_60_clock = clock;
  assign FF_60_reset = reset;
  assign FF_61_io_in = io_dram_wdata_bits_wdata_4;
  assign FF_61_io_init = 32'h5d6fc1;
  assign FF_61_io_enable = _T_1534;
  assign FF_61_clock = clock;
  assign FF_61_reset = reset;
  assign FF_62_io_in = io_dram_wdata_bits_wdata_5;
  assign FF_62_io_init = 32'h5d6fc2;
  assign FF_62_io_enable = _T_1534;
  assign FF_62_clock = clock;
  assign FF_62_reset = reset;
  assign FF_63_io_in = io_dram_wdata_bits_wdata_6;
  assign FF_63_io_init = 32'h5d6fc3;
  assign FF_63_io_enable = _T_1534;
  assign FF_63_clock = clock;
  assign FF_63_reset = reset;
  assign FF_64_io_in = io_dram_wdata_bits_wdata_7;
  assign FF_64_io_init = 32'h5d6fc4;
  assign FF_64_io_enable = _T_1534;
  assign FF_64_clock = clock;
  assign FF_64_reset = reset;
  assign FF_65_io_in = io_dram_wdata_bits_wdata_8;
  assign FF_65_io_init = 32'h5d6fc5;
  assign FF_65_io_enable = _T_1534;
  assign FF_65_clock = clock;
  assign FF_65_reset = reset;
  assign FF_66_io_in = io_dram_wdata_bits_wdata_9;
  assign FF_66_io_init = 32'h5d6fc6;
  assign FF_66_io_enable = _T_1534;
  assign FF_66_clock = clock;
  assign FF_66_reset = reset;
  assign FF_67_io_in = io_dram_wdata_bits_wdata_10;
  assign FF_67_io_init = 32'h5d6fc7;
  assign FF_67_io_enable = _T_1534;
  assign FF_67_clock = clock;
  assign FF_67_reset = reset;
  assign FF_68_io_in = io_dram_wdata_bits_wdata_11;
  assign FF_68_io_init = 32'h5d6fc8;
  assign FF_68_io_enable = _T_1534;
  assign FF_68_clock = clock;
  assign FF_68_reset = reset;
  assign FF_69_io_in = io_dram_wdata_bits_wdata_12;
  assign FF_69_io_init = 32'h5d6fc9;
  assign FF_69_io_enable = _T_1534;
  assign FF_69_clock = clock;
  assign FF_69_reset = reset;
  assign FF_70_io_in = io_dram_wdata_bits_wdata_13;
  assign FF_70_io_init = 32'h5d6fca;
  assign FF_70_io_enable = _T_1534;
  assign FF_70_clock = clock;
  assign FF_70_reset = reset;
  assign FF_71_io_in = io_dram_wdata_bits_wdata_14;
  assign FF_71_io_init = 32'h5d6fcb;
  assign FF_71_io_enable = _T_1534;
  assign FF_71_clock = clock;
  assign FF_71_reset = reset;
  assign FF_72_io_in = io_dram_wdata_bits_wdata_15;
  assign FF_72_io_init = 32'h5d6fcc;
  assign FF_72_io_enable = _T_1534;
  assign FF_72_clock = clock;
  assign FF_72_reset = reset;
  assign FF_73_io_in = _T_1527;
  assign FF_73_io_init = 512'h5d6fcd;
  assign FF_73_io_enable = _T_1534;
  assign FF_73_clock = clock;
  assign FF_73_reset = reset;
  assign Counter_3_io_max = 32'hffffffff;
  assign Counter_3_io_enable = _T_1666;
  assign Counter_3_clock = clock;
  assign Counter_3_reset = reset;
  assign Counter_4_io_max = 32'hffffffff;
  assign Counter_4_io_enable = _T_1676;
  assign Counter_4_clock = clock;
  assign Counter_4_reset = reset;
  assign Counter_5_io_max = 32'hffffffff;
  assign Counter_5_io_enable = _T_1685;
  assign Counter_5_clock = clock;
  assign Counter_5_reset = reset;
  assign Counter_6_io_max = 32'hffffffff;
  assign Counter_6_io_enable = 1'h0;
  assign Counter_6_clock = clock;
  assign Counter_6_reset = reset;
  assign Counter_7_io_max = 32'hffffffff;
  assign Counter_7_io_enable = 1'h0;
  assign Counter_7_clock = clock;
  assign Counter_7_reset = reset;
  assign Counter_8_io_max = 32'hffffffff;
  assign Counter_8_io_enable = _T_1707;
  assign Counter_8_clock = clock;
  assign Counter_8_reset = reset;
  assign Counter_9_io_max = 32'hffffffff;
  assign Counter_9_io_enable = _T_1715;
  assign Counter_9_clock = clock;
  assign Counter_9_reset = reset;
  assign Counter_10_io_max = 32'hffffffff;
  assign Counter_10_io_enable = 1'h0;
  assign Counter_10_clock = clock;
  assign Counter_10_reset = reset;
  assign Counter_11_io_max = 32'hffffffff;
  assign Counter_11_io_enable = 1'h0;
  assign Counter_11_clock = clock;
  assign Counter_11_reset = reset;
  assign Counter_12_io_max = 32'hffffffff;
  assign Counter_12_io_enable = _T_1737;
  assign Counter_12_clock = clock;
  assign Counter_12_reset = reset;
  assign Counter_13_io_max = 32'hffffffff;
  assign Counter_13_io_enable = _T_1160;
  assign Counter_13_clock = clock;
  assign Counter_13_reset = reset;
  assign Counter_14_io_max = 32'hffffffff;
  assign Counter_14_io_enable = _T_1751;
  assign Counter_14_clock = clock;
  assign Counter_14_reset = reset;
  assign Counter_15_io_max = 32'hffffffff;
  assign Counter_15_io_enable = _T_1759;
  assign Counter_15_clock = clock;
  assign Counter_15_reset = reset;
  assign Counter_16_io_max = 32'hffffffff;
  assign Counter_16_io_enable = _T_1768;
  assign Counter_16_clock = clock;
  assign Counter_16_reset = reset;
  assign Counter_17_io_max = 32'hffffffff;
  assign Counter_17_io_enable = _T_1774;
  assign Counter_17_clock = clock;
  assign Counter_17_reset = reset;
  assign Counter_18_io_max = 32'hffffffff;
  assign Counter_18_io_enable = _T_1782;
  assign Counter_18_clock = clock;
  assign Counter_18_reset = reset;
  assign Counter_19_io_max = 32'hffffffff;
  assign Counter_19_io_enable = _T_1790;
  assign Counter_19_clock = clock;
  assign Counter_19_reset = reset;
  assign Counter_20_io_max = 32'hffffffff;
  assign Counter_20_io_enable = _T_1799;
  assign Counter_20_clock = clock;
  assign Counter_20_reset = reset;
  assign Counter_21_io_max = 32'hffffffff;
  assign Counter_21_io_enable = denseLoadBuffers_0_io_full;
  assign Counter_21_clock = clock;
  assign Counter_21_reset = reset;
  assign Counter_22_io_max = 32'hffffffff;
  assign Counter_22_io_enable = denseLoadBuffers_0_io_almostFull;
  assign Counter_22_clock = clock;
  assign Counter_22_reset = reset;
  assign Counter_23_io_max = 32'hffffffff;
  assign Counter_23_io_enable = denseLoadBuffers_0_io_empty;
  assign Counter_23_clock = clock;
  assign Counter_23_reset = reset;
  assign Counter_24_io_max = 32'hffffffff;
  assign Counter_24_io_enable = denseLoadBuffers_0_io_almostEmpty;
  assign Counter_24_clock = clock;
  assign Counter_24_reset = reset;
  assign Counter_25_io_max = 32'hffffffff;
  assign Counter_25_io_enable = denseLoadBuffers_0_io_enqVld;
  assign Counter_25_clock = clock;
  assign Counter_25_reset = reset;
  assign Counter_26_io_max = 32'hffffffff;
  assign Counter_26_io_enable = _T_1035;
  assign Counter_26_clock = clock;
  assign Counter_26_reset = reset;
  assign Counter_27_io_max = 32'hffffffff;
  assign Counter_27_io_enable = io_dram_rresp_valid;
  assign Counter_27_clock = clock;
  assign Counter_27_reset = reset;
  assign Counter_28_io_max = 32'hffffffff;
  assign Counter_28_io_enable = _T_1843;
  assign Counter_28_clock = clock;
  assign Counter_28_reset = reset;
  assign FF_74_io_in = io_dram_rresp_bits_tag_streamId;
  assign FF_74_io_init = 6'h28;
  assign FF_74_io_enable = io_dram_rresp_valid;
  assign FF_74_clock = clock;
  assign FF_74_reset = reset;
  assign Counter_29_io_max = 32'hffffffff;
  assign Counter_29_io_enable = denseStoreBuffers_0_io_full;
  assign Counter_29_clock = clock;
  assign Counter_29_reset = reset;
  assign Counter_30_io_max = 32'hffffffff;
  assign Counter_30_io_enable = denseStoreBuffers_0_io_almostFull;
  assign Counter_30_clock = clock;
  assign Counter_30_reset = reset;
  assign Counter_31_io_max = 32'hffffffff;
  assign Counter_31_io_enable = denseStoreBuffers_0_io_empty;
  assign Counter_31_clock = clock;
  assign Counter_31_reset = reset;
  assign Counter_32_io_max = 32'hffffffff;
  assign Counter_32_io_enable = denseStoreBuffers_0_io_almostEmpty;
  assign Counter_32_clock = clock;
  assign Counter_32_reset = reset;
  assign Counter_33_io_max = 32'hffffffff;
  assign Counter_33_io_enable = _T_1872;
  assign Counter_33_clock = clock;
  assign Counter_33_reset = reset;
  assign Counter_34_io_max = 32'hffffffff;
  assign Counter_34_io_enable = _T_1160;
  assign Counter_34_clock = clock;
  assign Counter_34_reset = reset;
  assign Counter_35_io_max = 32'hffffffff;
  assign Counter_35_io_enable = _T_1885;
  assign Counter_35_clock = clock;
  assign Counter_35_reset = reset;
  assign Counter_36_io_max = 32'hffffffff;
  assign Counter_36_io_enable = _T_1892;
  assign Counter_36_clock = clock;
  assign Counter_36_reset = reset;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_1058 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_1088 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1058 <= 1'h0;
    end else begin
      _T_1058 <= _T_1055;
    end
    if (reset) begin
      _T_1088 <= 1'h0;
    end else begin
      _T_1088 <= _T_1085;
    end
  end
endmodule
module MuxN_16(
  input  [63:0] io_ins_0,
  input  [63:0] io_ins_1,
  input  [63:0] io_ins_2,
  input  [63:0] io_ins_3,
  input  [63:0] io_ins_4,
  input  [63:0] io_ins_5,
  input  [63:0] io_ins_6,
  input  [63:0] io_ins_7,
  input  [63:0] io_ins_8,
  input  [63:0] io_ins_9,
  input  [63:0] io_ins_10,
  input  [63:0] io_ins_11,
  input  [63:0] io_ins_12,
  input  [63:0] io_ins_13,
  input  [63:0] io_ins_14,
  input  [63:0] io_ins_15,
  input  [63:0] io_ins_16,
  input  [63:0] io_ins_17,
  input  [63:0] io_ins_18,
  input  [63:0] io_ins_19,
  input  [63:0] io_ins_20,
  input  [63:0] io_ins_21,
  input  [63:0] io_ins_22,
  input  [63:0] io_ins_23,
  input  [63:0] io_ins_24,
  input  [63:0] io_ins_25,
  input  [63:0] io_ins_26,
  input  [63:0] io_ins_27,
  input  [63:0] io_ins_28,
  input  [63:0] io_ins_29,
  input  [63:0] io_ins_30,
  input  [63:0] io_ins_31,
  input  [63:0] io_ins_32,
  input  [63:0] io_ins_33,
  input  [63:0] io_ins_34,
  input  [63:0] io_ins_35,
  input  [63:0] io_ins_36,
  input  [63:0] io_ins_37,
  input  [63:0] io_ins_38,
  input  [63:0] io_ins_39,
  input  [63:0] io_ins_40,
  input  [63:0] io_ins_41,
  input  [63:0] io_ins_42,
  input  [63:0] io_ins_43,
  input  [63:0] io_ins_44,
  input  [63:0] io_ins_45,
  input  [63:0] io_ins_46,
  input  [63:0] io_ins_47,
  input  [63:0] io_ins_48,
  input  [63:0] io_ins_49,
  input  [63:0] io_ins_50,
  input  [63:0] io_ins_51,
  input  [63:0] io_ins_52,
  input  [63:0] io_ins_53,
  input  [63:0] io_ins_54,
  input  [63:0] io_ins_55,
  input  [63:0] io_ins_56,
  input  [63:0] io_ins_57,
  input  [63:0] io_ins_58,
  input  [63:0] io_ins_59,
  input  [63:0] io_ins_60,
  input  [63:0] io_ins_61,
  input  [63:0] io_ins_62,
  input  [63:0] io_ins_63,
  input  [63:0] io_ins_64,
  input  [63:0] io_ins_65,
  input  [63:0] io_ins_66,
  input  [63:0] io_ins_67,
  input  [63:0] io_ins_68,
  input  [63:0] io_ins_69,
  input  [63:0] io_ins_70,
  input  [63:0] io_ins_71,
  input  [63:0] io_ins_72,
  input  [63:0] io_ins_73,
  input  [63:0] io_ins_74,
  input  [63:0] io_ins_75,
  input  [63:0] io_ins_76,
  input  [63:0] io_ins_77,
  input  [63:0] io_ins_78,
  input  [63:0] io_ins_79,
  input  [63:0] io_ins_80,
  input  [63:0] io_ins_81,
  input  [63:0] io_ins_82,
  input  [63:0] io_ins_83,
  input  [63:0] io_ins_84,
  input  [63:0] io_ins_85,
  input  [63:0] io_ins_86,
  input  [63:0] io_ins_87,
  input  [63:0] io_ins_88,
  input  [63:0] io_ins_89,
  input  [63:0] io_ins_90,
  input  [63:0] io_ins_91,
  input  [63:0] io_ins_92,
  input  [63:0] io_ins_93,
  input  [63:0] io_ins_94,
  input  [63:0] io_ins_95,
  input  [63:0] io_ins_96,
  input  [63:0] io_ins_97,
  input  [63:0] io_ins_98,
  input  [63:0] io_ins_99,
  input  [63:0] io_ins_100,
  input  [63:0] io_ins_101,
  input  [63:0] io_ins_102,
  input  [63:0] io_ins_103,
  input  [63:0] io_ins_104,
  input  [63:0] io_ins_105,
  input  [63:0] io_ins_106,
  input  [63:0] io_ins_107,
  input  [63:0] io_ins_108,
  input  [63:0] io_ins_109,
  input  [63:0] io_ins_110,
  input  [63:0] io_ins_111,
  input  [63:0] io_ins_112,
  input  [63:0] io_ins_113,
  input  [63:0] io_ins_114,
  input  [63:0] io_ins_115,
  input  [63:0] io_ins_116,
  input  [63:0] io_ins_117,
  input  [63:0] io_ins_118,
  input  [63:0] io_ins_119,
  input  [63:0] io_ins_120,
  input  [63:0] io_ins_121,
  input  [63:0] io_ins_122,
  input  [63:0] io_ins_123,
  input  [63:0] io_ins_124,
  input  [63:0] io_ins_125,
  input  [63:0] io_ins_126,
  input  [63:0] io_ins_127,
  input  [63:0] io_ins_128,
  input  [63:0] io_ins_129,
  input  [63:0] io_ins_130,
  input  [63:0] io_ins_131,
  input  [63:0] io_ins_132,
  input  [63:0] io_ins_133,
  input  [63:0] io_ins_134,
  input  [63:0] io_ins_135,
  input  [63:0] io_ins_136,
  input  [63:0] io_ins_137,
  input  [63:0] io_ins_138,
  input  [63:0] io_ins_139,
  input  [63:0] io_ins_140,
  input  [63:0] io_ins_141,
  input  [63:0] io_ins_142,
  input  [63:0] io_ins_143,
  input  [63:0] io_ins_144,
  input  [63:0] io_ins_145,
  input  [63:0] io_ins_146,
  input  [63:0] io_ins_147,
  input  [63:0] io_ins_148,
  input  [63:0] io_ins_149,
  input  [63:0] io_ins_150,
  input  [63:0] io_ins_151,
  input  [63:0] io_ins_152,
  input  [63:0] io_ins_153,
  input  [63:0] io_ins_154,
  input  [63:0] io_ins_155,
  input  [63:0] io_ins_156,
  input  [63:0] io_ins_157,
  input  [63:0] io_ins_158,
  input  [63:0] io_ins_159,
  input  [63:0] io_ins_160,
  input  [63:0] io_ins_161,
  input  [63:0] io_ins_162,
  input  [63:0] io_ins_163,
  input  [63:0] io_ins_164,
  input  [63:0] io_ins_165,
  input  [63:0] io_ins_166,
  input  [63:0] io_ins_167,
  input  [63:0] io_ins_168,
  input  [63:0] io_ins_169,
  input  [63:0] io_ins_170,
  input  [63:0] io_ins_171,
  input  [63:0] io_ins_172,
  input  [63:0] io_ins_173,
  input  [63:0] io_ins_174,
  input  [63:0] io_ins_175,
  input  [63:0] io_ins_176,
  input  [63:0] io_ins_177,
  input  [63:0] io_ins_178,
  input  [63:0] io_ins_179,
  input  [63:0] io_ins_180,
  input  [63:0] io_ins_181,
  input  [63:0] io_ins_182,
  input  [63:0] io_ins_183,
  input  [63:0] io_ins_184,
  input  [63:0] io_ins_185,
  input  [63:0] io_ins_186,
  input  [63:0] io_ins_187,
  input  [63:0] io_ins_188,
  input  [63:0] io_ins_189,
  input  [63:0] io_ins_190,
  input  [63:0] io_ins_191,
  input  [63:0] io_ins_192,
  input  [63:0] io_ins_193,
  input  [63:0] io_ins_194,
  input  [63:0] io_ins_195,
  input  [63:0] io_ins_196,
  input  [63:0] io_ins_197,
  input  [63:0] io_ins_198,
  input  [63:0] io_ins_199,
  input  [63:0] io_ins_200,
  input  [63:0] io_ins_201,
  input  [63:0] io_ins_202,
  input  [63:0] io_ins_203,
  input  [63:0] io_ins_204,
  input  [63:0] io_ins_205,
  input  [63:0] io_ins_206,
  input  [63:0] io_ins_207,
  input  [63:0] io_ins_208,
  input  [63:0] io_ins_209,
  input  [63:0] io_ins_210,
  input  [63:0] io_ins_211,
  input  [63:0] io_ins_212,
  input  [63:0] io_ins_213,
  input  [63:0] io_ins_214,
  input  [63:0] io_ins_215,
  input  [63:0] io_ins_216,
  input  [63:0] io_ins_217,
  input  [63:0] io_ins_218,
  input  [63:0] io_ins_219,
  input  [63:0] io_ins_220,
  input  [63:0] io_ins_221,
  input  [63:0] io_ins_222,
  input  [63:0] io_ins_223,
  input  [63:0] io_ins_224,
  input  [63:0] io_ins_225,
  input  [63:0] io_ins_226,
  input  [63:0] io_ins_227,
  input  [63:0] io_ins_228,
  input  [63:0] io_ins_229,
  input  [63:0] io_ins_230,
  input  [63:0] io_ins_231,
  input  [63:0] io_ins_232,
  input  [63:0] io_ins_233,
  input  [63:0] io_ins_234,
  input  [63:0] io_ins_235,
  input  [63:0] io_ins_236,
  input  [63:0] io_ins_237,
  input  [63:0] io_ins_238,
  input  [63:0] io_ins_239,
  input  [63:0] io_ins_240,
  input  [63:0] io_ins_241,
  input  [63:0] io_ins_242,
  input  [63:0] io_ins_243,
  input  [63:0] io_ins_244,
  input  [63:0] io_ins_245,
  input  [63:0] io_ins_246,
  input  [63:0] io_ins_247,
  input  [63:0] io_ins_248,
  input  [63:0] io_ins_249,
  input  [63:0] io_ins_250,
  input  [63:0] io_ins_251,
  input  [63:0] io_ins_252,
  input  [63:0] io_ins_253,
  input  [63:0] io_ins_254,
  input  [63:0] io_ins_255,
  input  [63:0] io_ins_256,
  input  [63:0] io_ins_257,
  input  [63:0] io_ins_258,
  input  [63:0] io_ins_259,
  input  [63:0] io_ins_260,
  input  [63:0] io_ins_261,
  input  [63:0] io_ins_262,
  input  [63:0] io_ins_263,
  input  [63:0] io_ins_264,
  input  [63:0] io_ins_265,
  input  [63:0] io_ins_266,
  input  [63:0] io_ins_267,
  input  [63:0] io_ins_268,
  input  [63:0] io_ins_269,
  input  [63:0] io_ins_270,
  input  [63:0] io_ins_271,
  input  [63:0] io_ins_272,
  input  [63:0] io_ins_273,
  input  [63:0] io_ins_274,
  input  [63:0] io_ins_275,
  input  [63:0] io_ins_276,
  input  [63:0] io_ins_277,
  input  [63:0] io_ins_278,
  input  [63:0] io_ins_279,
  input  [63:0] io_ins_280,
  input  [63:0] io_ins_281,
  input  [63:0] io_ins_282,
  input  [63:0] io_ins_283,
  input  [63:0] io_ins_284,
  input  [63:0] io_ins_285,
  input  [63:0] io_ins_286,
  input  [63:0] io_ins_287,
  input  [63:0] io_ins_288,
  input  [63:0] io_ins_289,
  input  [63:0] io_ins_290,
  input  [63:0] io_ins_291,
  input  [63:0] io_ins_292,
  input  [63:0] io_ins_293,
  input  [63:0] io_ins_294,
  input  [63:0] io_ins_295,
  input  [63:0] io_ins_296,
  input  [63:0] io_ins_297,
  input  [63:0] io_ins_298,
  input  [63:0] io_ins_299,
  input  [63:0] io_ins_300,
  input  [63:0] io_ins_301,
  input  [63:0] io_ins_302,
  input  [63:0] io_ins_303,
  input  [63:0] io_ins_304,
  input  [63:0] io_ins_305,
  input  [63:0] io_ins_306,
  input  [63:0] io_ins_307,
  input  [63:0] io_ins_308,
  input  [63:0] io_ins_309,
  input  [63:0] io_ins_310,
  input  [63:0] io_ins_311,
  input  [63:0] io_ins_312,
  input  [63:0] io_ins_313,
  input  [63:0] io_ins_314,
  input  [63:0] io_ins_315,
  input  [63:0] io_ins_316,
  input  [63:0] io_ins_317,
  input  [63:0] io_ins_318,
  input  [63:0] io_ins_319,
  input  [63:0] io_ins_320,
  input  [63:0] io_ins_321,
  input  [63:0] io_ins_322,
  input  [63:0] io_ins_323,
  input  [63:0] io_ins_324,
  input  [63:0] io_ins_325,
  input  [63:0] io_ins_326,
  input  [63:0] io_ins_327,
  input  [63:0] io_ins_328,
  input  [63:0] io_ins_329,
  input  [63:0] io_ins_330,
  input  [63:0] io_ins_331,
  input  [63:0] io_ins_332,
  input  [63:0] io_ins_333,
  input  [63:0] io_ins_334,
  input  [63:0] io_ins_335,
  input  [63:0] io_ins_336,
  input  [63:0] io_ins_337,
  input  [63:0] io_ins_338,
  input  [63:0] io_ins_339,
  input  [63:0] io_ins_340,
  input  [63:0] io_ins_341,
  input  [63:0] io_ins_342,
  input  [63:0] io_ins_343,
  input  [63:0] io_ins_344,
  input  [63:0] io_ins_345,
  input  [63:0] io_ins_346,
  input  [63:0] io_ins_347,
  input  [63:0] io_ins_348,
  input  [63:0] io_ins_349,
  input  [63:0] io_ins_350,
  input  [63:0] io_ins_351,
  input  [63:0] io_ins_352,
  input  [63:0] io_ins_353,
  input  [63:0] io_ins_354,
  input  [63:0] io_ins_355,
  input  [63:0] io_ins_356,
  input  [63:0] io_ins_357,
  input  [63:0] io_ins_358,
  input  [63:0] io_ins_359,
  input  [63:0] io_ins_360,
  input  [63:0] io_ins_361,
  input  [63:0] io_ins_362,
  input  [63:0] io_ins_363,
  input  [63:0] io_ins_364,
  input  [63:0] io_ins_365,
  input  [63:0] io_ins_366,
  input  [63:0] io_ins_367,
  input  [63:0] io_ins_368,
  input  [63:0] io_ins_369,
  input  [63:0] io_ins_370,
  input  [63:0] io_ins_371,
  input  [63:0] io_ins_372,
  input  [63:0] io_ins_373,
  input  [63:0] io_ins_374,
  input  [63:0] io_ins_375,
  input  [63:0] io_ins_376,
  input  [63:0] io_ins_377,
  input  [63:0] io_ins_378,
  input  [63:0] io_ins_379,
  input  [63:0] io_ins_380,
  input  [63:0] io_ins_381,
  input  [63:0] io_ins_382,
  input  [63:0] io_ins_383,
  input  [63:0] io_ins_384,
  input  [63:0] io_ins_385,
  input  [63:0] io_ins_386,
  input  [63:0] io_ins_387,
  input  [63:0] io_ins_388,
  input  [63:0] io_ins_389,
  input  [63:0] io_ins_390,
  input  [63:0] io_ins_391,
  input  [63:0] io_ins_392,
  input  [63:0] io_ins_393,
  input  [63:0] io_ins_394,
  input  [63:0] io_ins_395,
  input  [63:0] io_ins_396,
  input  [63:0] io_ins_397,
  input  [63:0] io_ins_398,
  input  [63:0] io_ins_399,
  input  [63:0] io_ins_400,
  input  [63:0] io_ins_401,
  input  [63:0] io_ins_402,
  input  [63:0] io_ins_403,
  input  [63:0] io_ins_404,
  input  [63:0] io_ins_405,
  input  [63:0] io_ins_406,
  input  [63:0] io_ins_407,
  input  [63:0] io_ins_408,
  input  [63:0] io_ins_409,
  input  [63:0] io_ins_410,
  input  [63:0] io_ins_411,
  input  [63:0] io_ins_412,
  input  [63:0] io_ins_413,
  input  [63:0] io_ins_414,
  input  [63:0] io_ins_415,
  input  [63:0] io_ins_416,
  input  [63:0] io_ins_417,
  input  [63:0] io_ins_418,
  input  [63:0] io_ins_419,
  input  [63:0] io_ins_420,
  input  [63:0] io_ins_421,
  input  [63:0] io_ins_422,
  input  [63:0] io_ins_423,
  input  [63:0] io_ins_424,
  input  [63:0] io_ins_425,
  input  [63:0] io_ins_426,
  input  [63:0] io_ins_427,
  input  [63:0] io_ins_428,
  input  [63:0] io_ins_429,
  input  [63:0] io_ins_430,
  input  [63:0] io_ins_431,
  input  [63:0] io_ins_432,
  input  [63:0] io_ins_433,
  input  [63:0] io_ins_434,
  input  [63:0] io_ins_435,
  input  [63:0] io_ins_436,
  input  [63:0] io_ins_437,
  input  [63:0] io_ins_438,
  input  [63:0] io_ins_439,
  input  [63:0] io_ins_440,
  input  [63:0] io_ins_441,
  input  [63:0] io_ins_442,
  input  [63:0] io_ins_443,
  input  [63:0] io_ins_444,
  input  [63:0] io_ins_445,
  input  [63:0] io_ins_446,
  input  [63:0] io_ins_447,
  input  [63:0] io_ins_448,
  input  [63:0] io_ins_449,
  input  [63:0] io_ins_450,
  input  [63:0] io_ins_451,
  input  [63:0] io_ins_452,
  input  [63:0] io_ins_453,
  input  [63:0] io_ins_454,
  input  [63:0] io_ins_455,
  input  [63:0] io_ins_456,
  input  [63:0] io_ins_457,
  input  [63:0] io_ins_458,
  input  [63:0] io_ins_459,
  input  [63:0] io_ins_460,
  input  [63:0] io_ins_461,
  input  [63:0] io_ins_462,
  input  [63:0] io_ins_463,
  input  [63:0] io_ins_464,
  input  [63:0] io_ins_465,
  input  [63:0] io_ins_466,
  input  [63:0] io_ins_467,
  input  [63:0] io_ins_468,
  input  [63:0] io_ins_469,
  input  [63:0] io_ins_470,
  input  [63:0] io_ins_471,
  input  [63:0] io_ins_472,
  input  [63:0] io_ins_473,
  input  [63:0] io_ins_474,
  input  [63:0] io_ins_475,
  input  [63:0] io_ins_476,
  input  [63:0] io_ins_477,
  input  [63:0] io_ins_478,
  input  [63:0] io_ins_479,
  input  [63:0] io_ins_480,
  input  [63:0] io_ins_481,
  input  [63:0] io_ins_482,
  input  [63:0] io_ins_483,
  input  [63:0] io_ins_484,
  input  [63:0] io_ins_485,
  input  [63:0] io_ins_486,
  input  [63:0] io_ins_487,
  input  [63:0] io_ins_488,
  input  [63:0] io_ins_489,
  input  [63:0] io_ins_490,
  input  [63:0] io_ins_491,
  input  [63:0] io_ins_492,
  input  [63:0] io_ins_493,
  input  [63:0] io_ins_494,
  input  [63:0] io_ins_495,
  input  [63:0] io_ins_496,
  input  [63:0] io_ins_497,
  input  [63:0] io_ins_498,
  input  [63:0] io_ins_499,
  input  [63:0] io_ins_500,
  input  [63:0] io_ins_501,
  input  [63:0] io_ins_502,
  input  [63:0] io_ins_503,
  input  [63:0] io_ins_504,
  input  [8:0]  io_sel,
  output [63:0] io_out
);
  wire [63:0] _GEN_0;
  wire [63:0] _GEN_1;
  wire [63:0] _GEN_2;
  wire [63:0] _GEN_3;
  wire [63:0] _GEN_4;
  wire [63:0] _GEN_5;
  wire [63:0] _GEN_6;
  wire [63:0] _GEN_7;
  wire [63:0] _GEN_8;
  wire [63:0] _GEN_9;
  wire [63:0] _GEN_10;
  wire [63:0] _GEN_11;
  wire [63:0] _GEN_12;
  wire [63:0] _GEN_13;
  wire [63:0] _GEN_14;
  wire [63:0] _GEN_15;
  wire [63:0] _GEN_16;
  wire [63:0] _GEN_17;
  wire [63:0] _GEN_18;
  wire [63:0] _GEN_19;
  wire [63:0] _GEN_20;
  wire [63:0] _GEN_21;
  wire [63:0] _GEN_22;
  wire [63:0] _GEN_23;
  wire [63:0] _GEN_24;
  wire [63:0] _GEN_25;
  wire [63:0] _GEN_26;
  wire [63:0] _GEN_27;
  wire [63:0] _GEN_28;
  wire [63:0] _GEN_29;
  wire [63:0] _GEN_30;
  wire [63:0] _GEN_31;
  wire [63:0] _GEN_32;
  wire [63:0] _GEN_33;
  wire [63:0] _GEN_34;
  wire [63:0] _GEN_35;
  wire [63:0] _GEN_36;
  wire [63:0] _GEN_37;
  wire [63:0] _GEN_38;
  wire [63:0] _GEN_39;
  wire [63:0] _GEN_40;
  wire [63:0] _GEN_41;
  wire [63:0] _GEN_42;
  wire [63:0] _GEN_43;
  wire [63:0] _GEN_44;
  wire [63:0] _GEN_45;
  wire [63:0] _GEN_46;
  wire [63:0] _GEN_47;
  wire [63:0] _GEN_48;
  wire [63:0] _GEN_49;
  wire [63:0] _GEN_50;
  wire [63:0] _GEN_51;
  wire [63:0] _GEN_52;
  wire [63:0] _GEN_53;
  wire [63:0] _GEN_54;
  wire [63:0] _GEN_55;
  wire [63:0] _GEN_56;
  wire [63:0] _GEN_57;
  wire [63:0] _GEN_58;
  wire [63:0] _GEN_59;
  wire [63:0] _GEN_60;
  wire [63:0] _GEN_61;
  wire [63:0] _GEN_62;
  wire [63:0] _GEN_63;
  wire [63:0] _GEN_64;
  wire [63:0] _GEN_65;
  wire [63:0] _GEN_66;
  wire [63:0] _GEN_67;
  wire [63:0] _GEN_68;
  wire [63:0] _GEN_69;
  wire [63:0] _GEN_70;
  wire [63:0] _GEN_71;
  wire [63:0] _GEN_72;
  wire [63:0] _GEN_73;
  wire [63:0] _GEN_74;
  wire [63:0] _GEN_75;
  wire [63:0] _GEN_76;
  wire [63:0] _GEN_77;
  wire [63:0] _GEN_78;
  wire [63:0] _GEN_79;
  wire [63:0] _GEN_80;
  wire [63:0] _GEN_81;
  wire [63:0] _GEN_82;
  wire [63:0] _GEN_83;
  wire [63:0] _GEN_84;
  wire [63:0] _GEN_85;
  wire [63:0] _GEN_86;
  wire [63:0] _GEN_87;
  wire [63:0] _GEN_88;
  wire [63:0] _GEN_89;
  wire [63:0] _GEN_90;
  wire [63:0] _GEN_91;
  wire [63:0] _GEN_92;
  wire [63:0] _GEN_93;
  wire [63:0] _GEN_94;
  wire [63:0] _GEN_95;
  wire [63:0] _GEN_96;
  wire [63:0] _GEN_97;
  wire [63:0] _GEN_98;
  wire [63:0] _GEN_99;
  wire [63:0] _GEN_100;
  wire [63:0] _GEN_101;
  wire [63:0] _GEN_102;
  wire [63:0] _GEN_103;
  wire [63:0] _GEN_104;
  wire [63:0] _GEN_105;
  wire [63:0] _GEN_106;
  wire [63:0] _GEN_107;
  wire [63:0] _GEN_108;
  wire [63:0] _GEN_109;
  wire [63:0] _GEN_110;
  wire [63:0] _GEN_111;
  wire [63:0] _GEN_112;
  wire [63:0] _GEN_113;
  wire [63:0] _GEN_114;
  wire [63:0] _GEN_115;
  wire [63:0] _GEN_116;
  wire [63:0] _GEN_117;
  wire [63:0] _GEN_118;
  wire [63:0] _GEN_119;
  wire [63:0] _GEN_120;
  wire [63:0] _GEN_121;
  wire [63:0] _GEN_122;
  wire [63:0] _GEN_123;
  wire [63:0] _GEN_124;
  wire [63:0] _GEN_125;
  wire [63:0] _GEN_126;
  wire [63:0] _GEN_127;
  wire [63:0] _GEN_128;
  wire [63:0] _GEN_129;
  wire [63:0] _GEN_130;
  wire [63:0] _GEN_131;
  wire [63:0] _GEN_132;
  wire [63:0] _GEN_133;
  wire [63:0] _GEN_134;
  wire [63:0] _GEN_135;
  wire [63:0] _GEN_136;
  wire [63:0] _GEN_137;
  wire [63:0] _GEN_138;
  wire [63:0] _GEN_139;
  wire [63:0] _GEN_140;
  wire [63:0] _GEN_141;
  wire [63:0] _GEN_142;
  wire [63:0] _GEN_143;
  wire [63:0] _GEN_144;
  wire [63:0] _GEN_145;
  wire [63:0] _GEN_146;
  wire [63:0] _GEN_147;
  wire [63:0] _GEN_148;
  wire [63:0] _GEN_149;
  wire [63:0] _GEN_150;
  wire [63:0] _GEN_151;
  wire [63:0] _GEN_152;
  wire [63:0] _GEN_153;
  wire [63:0] _GEN_154;
  wire [63:0] _GEN_155;
  wire [63:0] _GEN_156;
  wire [63:0] _GEN_157;
  wire [63:0] _GEN_158;
  wire [63:0] _GEN_159;
  wire [63:0] _GEN_160;
  wire [63:0] _GEN_161;
  wire [63:0] _GEN_162;
  wire [63:0] _GEN_163;
  wire [63:0] _GEN_164;
  wire [63:0] _GEN_165;
  wire [63:0] _GEN_166;
  wire [63:0] _GEN_167;
  wire [63:0] _GEN_168;
  wire [63:0] _GEN_169;
  wire [63:0] _GEN_170;
  wire [63:0] _GEN_171;
  wire [63:0] _GEN_172;
  wire [63:0] _GEN_173;
  wire [63:0] _GEN_174;
  wire [63:0] _GEN_175;
  wire [63:0] _GEN_176;
  wire [63:0] _GEN_177;
  wire [63:0] _GEN_178;
  wire [63:0] _GEN_179;
  wire [63:0] _GEN_180;
  wire [63:0] _GEN_181;
  wire [63:0] _GEN_182;
  wire [63:0] _GEN_183;
  wire [63:0] _GEN_184;
  wire [63:0] _GEN_185;
  wire [63:0] _GEN_186;
  wire [63:0] _GEN_187;
  wire [63:0] _GEN_188;
  wire [63:0] _GEN_189;
  wire [63:0] _GEN_190;
  wire [63:0] _GEN_191;
  wire [63:0] _GEN_192;
  wire [63:0] _GEN_193;
  wire [63:0] _GEN_194;
  wire [63:0] _GEN_195;
  wire [63:0] _GEN_196;
  wire [63:0] _GEN_197;
  wire [63:0] _GEN_198;
  wire [63:0] _GEN_199;
  wire [63:0] _GEN_200;
  wire [63:0] _GEN_201;
  wire [63:0] _GEN_202;
  wire [63:0] _GEN_203;
  wire [63:0] _GEN_204;
  wire [63:0] _GEN_205;
  wire [63:0] _GEN_206;
  wire [63:0] _GEN_207;
  wire [63:0] _GEN_208;
  wire [63:0] _GEN_209;
  wire [63:0] _GEN_210;
  wire [63:0] _GEN_211;
  wire [63:0] _GEN_212;
  wire [63:0] _GEN_213;
  wire [63:0] _GEN_214;
  wire [63:0] _GEN_215;
  wire [63:0] _GEN_216;
  wire [63:0] _GEN_217;
  wire [63:0] _GEN_218;
  wire [63:0] _GEN_219;
  wire [63:0] _GEN_220;
  wire [63:0] _GEN_221;
  wire [63:0] _GEN_222;
  wire [63:0] _GEN_223;
  wire [63:0] _GEN_224;
  wire [63:0] _GEN_225;
  wire [63:0] _GEN_226;
  wire [63:0] _GEN_227;
  wire [63:0] _GEN_228;
  wire [63:0] _GEN_229;
  wire [63:0] _GEN_230;
  wire [63:0] _GEN_231;
  wire [63:0] _GEN_232;
  wire [63:0] _GEN_233;
  wire [63:0] _GEN_234;
  wire [63:0] _GEN_235;
  wire [63:0] _GEN_236;
  wire [63:0] _GEN_237;
  wire [63:0] _GEN_238;
  wire [63:0] _GEN_239;
  wire [63:0] _GEN_240;
  wire [63:0] _GEN_241;
  wire [63:0] _GEN_242;
  wire [63:0] _GEN_243;
  wire [63:0] _GEN_244;
  wire [63:0] _GEN_245;
  wire [63:0] _GEN_246;
  wire [63:0] _GEN_247;
  wire [63:0] _GEN_248;
  wire [63:0] _GEN_249;
  wire [63:0] _GEN_250;
  wire [63:0] _GEN_251;
  wire [63:0] _GEN_252;
  wire [63:0] _GEN_253;
  wire [63:0] _GEN_254;
  wire [63:0] _GEN_255;
  wire [63:0] _GEN_256;
  wire [63:0] _GEN_257;
  wire [63:0] _GEN_258;
  wire [63:0] _GEN_259;
  wire [63:0] _GEN_260;
  wire [63:0] _GEN_261;
  wire [63:0] _GEN_262;
  wire [63:0] _GEN_263;
  wire [63:0] _GEN_264;
  wire [63:0] _GEN_265;
  wire [63:0] _GEN_266;
  wire [63:0] _GEN_267;
  wire [63:0] _GEN_268;
  wire [63:0] _GEN_269;
  wire [63:0] _GEN_270;
  wire [63:0] _GEN_271;
  wire [63:0] _GEN_272;
  wire [63:0] _GEN_273;
  wire [63:0] _GEN_274;
  wire [63:0] _GEN_275;
  wire [63:0] _GEN_276;
  wire [63:0] _GEN_277;
  wire [63:0] _GEN_278;
  wire [63:0] _GEN_279;
  wire [63:0] _GEN_280;
  wire [63:0] _GEN_281;
  wire [63:0] _GEN_282;
  wire [63:0] _GEN_283;
  wire [63:0] _GEN_284;
  wire [63:0] _GEN_285;
  wire [63:0] _GEN_286;
  wire [63:0] _GEN_287;
  wire [63:0] _GEN_288;
  wire [63:0] _GEN_289;
  wire [63:0] _GEN_290;
  wire [63:0] _GEN_291;
  wire [63:0] _GEN_292;
  wire [63:0] _GEN_293;
  wire [63:0] _GEN_294;
  wire [63:0] _GEN_295;
  wire [63:0] _GEN_296;
  wire [63:0] _GEN_297;
  wire [63:0] _GEN_298;
  wire [63:0] _GEN_299;
  wire [63:0] _GEN_300;
  wire [63:0] _GEN_301;
  wire [63:0] _GEN_302;
  wire [63:0] _GEN_303;
  wire [63:0] _GEN_304;
  wire [63:0] _GEN_305;
  wire [63:0] _GEN_306;
  wire [63:0] _GEN_307;
  wire [63:0] _GEN_308;
  wire [63:0] _GEN_309;
  wire [63:0] _GEN_310;
  wire [63:0] _GEN_311;
  wire [63:0] _GEN_312;
  wire [63:0] _GEN_313;
  wire [63:0] _GEN_314;
  wire [63:0] _GEN_315;
  wire [63:0] _GEN_316;
  wire [63:0] _GEN_317;
  wire [63:0] _GEN_318;
  wire [63:0] _GEN_319;
  wire [63:0] _GEN_320;
  wire [63:0] _GEN_321;
  wire [63:0] _GEN_322;
  wire [63:0] _GEN_323;
  wire [63:0] _GEN_324;
  wire [63:0] _GEN_325;
  wire [63:0] _GEN_326;
  wire [63:0] _GEN_327;
  wire [63:0] _GEN_328;
  wire [63:0] _GEN_329;
  wire [63:0] _GEN_330;
  wire [63:0] _GEN_331;
  wire [63:0] _GEN_332;
  wire [63:0] _GEN_333;
  wire [63:0] _GEN_334;
  wire [63:0] _GEN_335;
  wire [63:0] _GEN_336;
  wire [63:0] _GEN_337;
  wire [63:0] _GEN_338;
  wire [63:0] _GEN_339;
  wire [63:0] _GEN_340;
  wire [63:0] _GEN_341;
  wire [63:0] _GEN_342;
  wire [63:0] _GEN_343;
  wire [63:0] _GEN_344;
  wire [63:0] _GEN_345;
  wire [63:0] _GEN_346;
  wire [63:0] _GEN_347;
  wire [63:0] _GEN_348;
  wire [63:0] _GEN_349;
  wire [63:0] _GEN_350;
  wire [63:0] _GEN_351;
  wire [63:0] _GEN_352;
  wire [63:0] _GEN_353;
  wire [63:0] _GEN_354;
  wire [63:0] _GEN_355;
  wire [63:0] _GEN_356;
  wire [63:0] _GEN_357;
  wire [63:0] _GEN_358;
  wire [63:0] _GEN_359;
  wire [63:0] _GEN_360;
  wire [63:0] _GEN_361;
  wire [63:0] _GEN_362;
  wire [63:0] _GEN_363;
  wire [63:0] _GEN_364;
  wire [63:0] _GEN_365;
  wire [63:0] _GEN_366;
  wire [63:0] _GEN_367;
  wire [63:0] _GEN_368;
  wire [63:0] _GEN_369;
  wire [63:0] _GEN_370;
  wire [63:0] _GEN_371;
  wire [63:0] _GEN_372;
  wire [63:0] _GEN_373;
  wire [63:0] _GEN_374;
  wire [63:0] _GEN_375;
  wire [63:0] _GEN_376;
  wire [63:0] _GEN_377;
  wire [63:0] _GEN_378;
  wire [63:0] _GEN_379;
  wire [63:0] _GEN_380;
  wire [63:0] _GEN_381;
  wire [63:0] _GEN_382;
  wire [63:0] _GEN_383;
  wire [63:0] _GEN_384;
  wire [63:0] _GEN_385;
  wire [63:0] _GEN_386;
  wire [63:0] _GEN_387;
  wire [63:0] _GEN_388;
  wire [63:0] _GEN_389;
  wire [63:0] _GEN_390;
  wire [63:0] _GEN_391;
  wire [63:0] _GEN_392;
  wire [63:0] _GEN_393;
  wire [63:0] _GEN_394;
  wire [63:0] _GEN_395;
  wire [63:0] _GEN_396;
  wire [63:0] _GEN_397;
  wire [63:0] _GEN_398;
  wire [63:0] _GEN_399;
  wire [63:0] _GEN_400;
  wire [63:0] _GEN_401;
  wire [63:0] _GEN_402;
  wire [63:0] _GEN_403;
  wire [63:0] _GEN_404;
  wire [63:0] _GEN_405;
  wire [63:0] _GEN_406;
  wire [63:0] _GEN_407;
  wire [63:0] _GEN_408;
  wire [63:0] _GEN_409;
  wire [63:0] _GEN_410;
  wire [63:0] _GEN_411;
  wire [63:0] _GEN_412;
  wire [63:0] _GEN_413;
  wire [63:0] _GEN_414;
  wire [63:0] _GEN_415;
  wire [63:0] _GEN_416;
  wire [63:0] _GEN_417;
  wire [63:0] _GEN_418;
  wire [63:0] _GEN_419;
  wire [63:0] _GEN_420;
  wire [63:0] _GEN_421;
  wire [63:0] _GEN_422;
  wire [63:0] _GEN_423;
  wire [63:0] _GEN_424;
  wire [63:0] _GEN_425;
  wire [63:0] _GEN_426;
  wire [63:0] _GEN_427;
  wire [63:0] _GEN_428;
  wire [63:0] _GEN_429;
  wire [63:0] _GEN_430;
  wire [63:0] _GEN_431;
  wire [63:0] _GEN_432;
  wire [63:0] _GEN_433;
  wire [63:0] _GEN_434;
  wire [63:0] _GEN_435;
  wire [63:0] _GEN_436;
  wire [63:0] _GEN_437;
  wire [63:0] _GEN_438;
  wire [63:0] _GEN_439;
  wire [63:0] _GEN_440;
  wire [63:0] _GEN_441;
  wire [63:0] _GEN_442;
  wire [63:0] _GEN_443;
  wire [63:0] _GEN_444;
  wire [63:0] _GEN_445;
  wire [63:0] _GEN_446;
  wire [63:0] _GEN_447;
  wire [63:0] _GEN_448;
  wire [63:0] _GEN_449;
  wire [63:0] _GEN_450;
  wire [63:0] _GEN_451;
  wire [63:0] _GEN_452;
  wire [63:0] _GEN_453;
  wire [63:0] _GEN_454;
  wire [63:0] _GEN_455;
  wire [63:0] _GEN_456;
  wire [63:0] _GEN_457;
  wire [63:0] _GEN_458;
  wire [63:0] _GEN_459;
  wire [63:0] _GEN_460;
  wire [63:0] _GEN_461;
  wire [63:0] _GEN_462;
  wire [63:0] _GEN_463;
  wire [63:0] _GEN_464;
  wire [63:0] _GEN_465;
  wire [63:0] _GEN_466;
  wire [63:0] _GEN_467;
  wire [63:0] _GEN_468;
  wire [63:0] _GEN_469;
  wire [63:0] _GEN_470;
  wire [63:0] _GEN_471;
  wire [63:0] _GEN_472;
  wire [63:0] _GEN_473;
  wire [63:0] _GEN_474;
  wire [63:0] _GEN_475;
  wire [63:0] _GEN_476;
  wire [63:0] _GEN_477;
  wire [63:0] _GEN_478;
  wire [63:0] _GEN_479;
  wire [63:0] _GEN_480;
  wire [63:0] _GEN_481;
  wire [63:0] _GEN_482;
  wire [63:0] _GEN_483;
  wire [63:0] _GEN_484;
  wire [63:0] _GEN_485;
  wire [63:0] _GEN_486;
  wire [63:0] _GEN_487;
  wire [63:0] _GEN_488;
  wire [63:0] _GEN_489;
  wire [63:0] _GEN_490;
  wire [63:0] _GEN_491;
  wire [63:0] _GEN_492;
  wire [63:0] _GEN_493;
  wire [63:0] _GEN_494;
  wire [63:0] _GEN_495;
  wire [63:0] _GEN_496;
  wire [63:0] _GEN_497;
  wire [63:0] _GEN_498;
  wire [63:0] _GEN_499;
  wire [63:0] _GEN_500;
  wire [63:0] _GEN_501;
  wire [63:0] _GEN_502;
  wire [63:0] _GEN_503;
  wire [63:0] _GEN_504;
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0;
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1;
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2;
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3;
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4;
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5;
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6;
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7;
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8;
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9;
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10;
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11;
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12;
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13;
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14;
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15;
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16;
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17;
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18;
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19;
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20;
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21;
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22;
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23;
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24;
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25;
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26;
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27;
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28;
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29;
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30;
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31;
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32;
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33;
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34;
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35;
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36;
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37;
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38;
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39;
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40;
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41;
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42;
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43;
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44;
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45;
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46;
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47;
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48;
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49;
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50;
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51;
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52;
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53;
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54;
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55;
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56;
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57;
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58;
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59;
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60;
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61;
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62;
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63;
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64;
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65;
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66;
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67;
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68;
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69;
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70;
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71;
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72;
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73;
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74;
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75;
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76;
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77;
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78;
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79;
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80;
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81;
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82;
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83;
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84;
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85;
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86;
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87;
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88;
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89;
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90;
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91;
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92;
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93;
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94;
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95;
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96;
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97;
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98;
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99;
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100;
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101;
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102;
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103;
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104;
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105;
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106;
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107;
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108;
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109;
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110;
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111;
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112;
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113;
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114;
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115;
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116;
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117;
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118;
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119;
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120;
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121;
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122;
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123;
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124;
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125;
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126;
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127;
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128;
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129;
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130;
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131;
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132;
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133;
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134;
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135;
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136;
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137;
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138;
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139;
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140;
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141;
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142;
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143;
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144;
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145;
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146;
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147;
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148;
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149;
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150;
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151;
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152;
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153;
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154;
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155;
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156;
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157;
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158;
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159;
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160;
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161;
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162;
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163;
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164;
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165;
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166;
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167;
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168;
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169;
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170;
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171;
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172;
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173;
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174;
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175;
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176;
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177;
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178;
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179;
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180;
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181;
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182;
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183;
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184;
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185;
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186;
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187;
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188;
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189;
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190;
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191;
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192;
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193;
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194;
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195;
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196;
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197;
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198;
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199;
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200;
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201;
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202;
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203;
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204;
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205;
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206;
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207;
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208;
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209;
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210;
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211;
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212;
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213;
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214;
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215;
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216;
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217;
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218;
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219;
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220;
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221;
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222;
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223;
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224;
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225;
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226;
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227;
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228;
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229;
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230;
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231;
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232;
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233;
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234;
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235;
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236;
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237;
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238;
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239;
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240;
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241;
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242;
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243;
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244;
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245;
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246;
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247;
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248;
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249;
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250;
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251;
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252;
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253;
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254;
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255;
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256;
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257;
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258;
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259;
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260;
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261;
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262;
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263;
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264;
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265;
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266;
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267;
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268;
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269;
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270;
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271;
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272;
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273;
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274;
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275;
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276;
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277;
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278;
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279;
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280;
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281;
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282;
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283;
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284;
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285;
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286;
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287;
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288;
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289;
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290;
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291;
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292;
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293;
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294;
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295;
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296;
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297;
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298;
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299;
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300;
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301;
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302;
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303;
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304;
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305;
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306;
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307;
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308;
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309;
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310;
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311;
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312;
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313;
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314;
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315;
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316;
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317;
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318;
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319;
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320;
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321;
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322;
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323;
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324;
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325;
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326;
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327;
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328;
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329;
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330;
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331;
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332;
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333;
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334;
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335;
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336;
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337;
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338;
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339;
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340;
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341;
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342;
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343;
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344;
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345;
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346;
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347;
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348;
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349;
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350;
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351;
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352;
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353;
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354;
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355;
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356;
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357;
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358;
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359;
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360;
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361;
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362;
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363;
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364;
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365;
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366;
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367;
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368;
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369;
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370;
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371;
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372;
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373;
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374;
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375;
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376;
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377;
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378;
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379;
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380;
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381;
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382;
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383;
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384;
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385;
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386;
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387;
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388;
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389;
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390;
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391;
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392;
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393;
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394;
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395;
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396;
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397;
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398;
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399;
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400;
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401;
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402;
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403;
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404;
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405;
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406;
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407;
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408;
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409;
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410;
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411;
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412;
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413;
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414;
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415;
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416;
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417;
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418;
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419;
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420;
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421;
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422;
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423;
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424;
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425;
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426;
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427;
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428;
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429;
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430;
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431;
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432;
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433;
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434;
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435;
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436;
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437;
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438;
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439;
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440;
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441;
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442;
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443;
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444;
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445;
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446;
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447;
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448;
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449;
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450;
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451;
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452;
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453;
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454;
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455;
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456;
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457;
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458;
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459;
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460;
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461;
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462;
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463;
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464;
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465;
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466;
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467;
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468;
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469;
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470;
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471;
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472;
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473;
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474;
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475;
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476;
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477;
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478;
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479;
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480;
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481;
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482;
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483;
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484;
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485;
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486;
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487;
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488;
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489;
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490;
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491;
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492;
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493;
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494;
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495;
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496;
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497;
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498;
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499;
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500;
  assign _GEN_502 = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501;
  assign _GEN_503 = 9'h1f7 == io_sel ? io_ins_503 : _GEN_502;
  assign _GEN_504 = 9'h1f8 == io_sel ? io_ins_504 : _GEN_503;
  assign io_out = _GEN_0;
  assign _GEN_0 = _GEN_504;
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [8:0]  io_raddr,
  input         io_wen,
  input  [8:0]  io_waddr,
  input  [63:0] io_wdata,
  output [63:0] io_rdata,
  output [63:0] io_argIns_0,
  output [63:0] io_argIns_1,
  output [63:0] io_argIns_2,
  output [63:0] io_argIns_3,
  input         io_argOuts_0_valid,
  input  [63:0] io_argOuts_0_bits,
  input         io_argOuts_1_valid,
  input  [63:0] io_argOuts_1_bits,
  input  [63:0] io_argOuts_2_bits,
  input  [63:0] io_argOuts_3_bits,
  input  [63:0] io_argOuts_4_bits,
  input  [63:0] io_argOuts_5_bits,
  input  [63:0] io_argOuts_6_bits,
  input  [63:0] io_argOuts_7_bits,
  input  [63:0] io_argOuts_8_bits,
  input  [63:0] io_argOuts_9_bits,
  input  [63:0] io_argOuts_10_bits,
  input  [63:0] io_argOuts_11_bits,
  input  [63:0] io_argOuts_12_bits,
  input  [63:0] io_argOuts_13_bits,
  input  [63:0] io_argOuts_14_bits,
  input  [63:0] io_argOuts_15_bits,
  input  [63:0] io_argOuts_16_bits,
  input  [63:0] io_argOuts_17_bits,
  input  [63:0] io_argOuts_18_bits,
  input  [63:0] io_argOuts_19_bits,
  input  [63:0] io_argOuts_20_bits,
  input  [63:0] io_argOuts_21_bits,
  input  [63:0] io_argOuts_22_bits,
  input  [63:0] io_argOuts_23_bits,
  input  [63:0] io_argOuts_24_bits,
  input  [63:0] io_argOuts_25_bits,
  input  [63:0] io_argOuts_26_bits,
  input  [63:0] io_argOuts_27_bits,
  input  [63:0] io_argOuts_28_bits,
  input  [63:0] io_argOuts_29_bits,
  input  [63:0] io_argOuts_30_bits,
  input  [63:0] io_argOuts_31_bits,
  input  [63:0] io_argOuts_32_bits,
  input  [63:0] io_argOuts_33_bits,
  input  [63:0] io_argOuts_34_bits,
  input  [63:0] io_argOuts_35_bits,
  input  [63:0] io_argOuts_36_bits,
  input  [63:0] io_argOuts_37_bits,
  input  [63:0] io_argOuts_38_bits,
  input  [63:0] io_argOuts_39_bits,
  input  [63:0] io_argOuts_40_bits,
  input  [63:0] io_argOuts_41_bits,
  input  [63:0] io_argOuts_42_bits,
  input  [63:0] io_argOuts_43_bits,
  input  [63:0] io_argOuts_44_bits,
  input  [63:0] io_argOuts_45_bits,
  input  [63:0] io_argOuts_46_bits,
  input  [63:0] io_argOuts_47_bits,
  input  [63:0] io_argOuts_48_bits,
  input  [63:0] io_argOuts_49_bits,
  input  [63:0] io_argOuts_50_bits,
  input  [63:0] io_argOuts_51_bits,
  input  [63:0] io_argOuts_52_bits,
  input  [63:0] io_argOuts_53_bits,
  input  [63:0] io_argOuts_54_bits,
  input  [63:0] io_argOuts_55_bits,
  input  [63:0] io_argOuts_56_bits,
  input  [63:0] io_argOuts_57_bits,
  input  [63:0] io_argOuts_58_bits,
  input  [63:0] io_argOuts_59_bits,
  input  [63:0] io_argOuts_60_bits,
  input  [63:0] io_argOuts_61_bits,
  input  [63:0] io_argOuts_62_bits,
  input  [63:0] io_argOuts_63_bits,
  input  [63:0] io_argOuts_64_bits,
  input  [63:0] io_argOuts_65_bits,
  input  [63:0] io_argOuts_66_bits,
  input  [63:0] io_argOuts_67_bits,
  input  [63:0] io_argOuts_68_bits,
  input  [63:0] io_argOuts_69_bits,
  input  [63:0] io_argOuts_70_bits,
  input  [63:0] io_argOuts_71_bits,
  input  [63:0] io_argOuts_72_bits,
  input  [63:0] io_argOuts_73_bits,
  input  [63:0] io_argOuts_74_bits,
  input  [63:0] io_argOuts_75_bits,
  input  [63:0] io_argOuts_76_bits,
  input  [63:0] io_argOuts_77_bits,
  input  [63:0] io_argOuts_78_bits,
  input  [63:0] io_argOuts_79_bits,
  input  [63:0] io_argOuts_80_bits,
  input  [63:0] io_argOuts_81_bits,
  input  [63:0] io_argOuts_82_bits,
  input  [63:0] io_argOuts_83_bits,
  input  [63:0] io_argOuts_84_bits,
  input  [63:0] io_argOuts_85_bits,
  input  [63:0] io_argOuts_86_bits,
  input  [63:0] io_argOuts_87_bits,
  input  [63:0] io_argOuts_88_bits,
  input  [63:0] io_argOuts_89_bits,
  input  [63:0] io_argOuts_90_bits,
  input  [63:0] io_argOuts_91_bits,
  input  [63:0] io_argOuts_92_bits,
  input  [63:0] io_argOuts_93_bits,
  input  [63:0] io_argOuts_94_bits,
  input  [63:0] io_argOuts_95_bits,
  input  [63:0] io_argOuts_96_bits,
  input  [63:0] io_argOuts_97_bits,
  input  [63:0] io_argOuts_98_bits,
  input  [63:0] io_argOuts_99_bits,
  input  [63:0] io_argOuts_100_bits,
  input  [63:0] io_argOuts_101_bits,
  input  [63:0] io_argOuts_102_bits,
  input  [63:0] io_argOuts_103_bits,
  input  [63:0] io_argOuts_104_bits,
  input  [63:0] io_argOuts_105_bits,
  input  [63:0] io_argOuts_106_bits,
  input  [63:0] io_argOuts_107_bits,
  input  [63:0] io_argOuts_108_bits,
  input  [63:0] io_argOuts_109_bits,
  input  [63:0] io_argOuts_110_bits,
  input  [63:0] io_argOuts_111_bits,
  input  [63:0] io_argOuts_112_bits,
  input  [63:0] io_argOuts_113_bits,
  input  [63:0] io_argOuts_114_bits,
  input  [63:0] io_argOuts_115_bits
);
  wire  regs_0_clock;
  wire  regs_0_reset;
  wire [63:0] regs_0_io_in;
  wire [63:0] regs_0_io_init;
  wire [63:0] regs_0_io_out;
  wire  regs_0_io_enable;
  wire  _T_1542;
  wire  _T_1543;
  wire  regs_1_clock;
  wire  regs_1_reset;
  wire [63:0] regs_1_io_in;
  wire [63:0] regs_1_io_init;
  wire [63:0] regs_1_io_out;
  wire  regs_1_io_enable;
  wire  _T_1546;
  wire  _T_1547;
  wire  _T_1551;
  wire [63:0] _T_1555;
  wire  regs_2_clock;
  wire  regs_2_reset;
  wire [63:0] regs_2_io_in;
  wire [63:0] regs_2_io_init;
  wire [63:0] regs_2_io_out;
  wire  regs_2_io_enable;
  wire  _T_1558;
  wire  _T_1559;
  wire  regs_3_clock;
  wire  regs_3_reset;
  wire [63:0] regs_3_io_in;
  wire [63:0] regs_3_io_init;
  wire [63:0] regs_3_io_out;
  wire  regs_3_io_enable;
  wire  _T_1562;
  wire  _T_1563;
  wire  regs_4_clock;
  wire  regs_4_reset;
  wire [63:0] regs_4_io_in;
  wire [63:0] regs_4_io_init;
  wire [63:0] regs_4_io_out;
  wire  regs_4_io_enable;
  wire  _T_1566;
  wire  _T_1567;
  wire  _T_1568;
  wire [63:0] _T_1569;
  wire  regs_5_clock;
  wire  regs_5_reset;
  wire [63:0] regs_5_io_in;
  wire [63:0] regs_5_io_init;
  wire [63:0] regs_5_io_out;
  wire  regs_5_io_enable;
  wire  regs_6_clock;
  wire  regs_6_reset;
  wire [63:0] regs_6_io_in;
  wire [63:0] regs_6_io_init;
  wire [63:0] regs_6_io_out;
  wire  regs_6_io_enable;
  wire  regs_7_clock;
  wire  regs_7_reset;
  wire [63:0] regs_7_io_in;
  wire [63:0] regs_7_io_init;
  wire [63:0] regs_7_io_out;
  wire  regs_7_io_enable;
  wire  regs_8_clock;
  wire  regs_8_reset;
  wire [63:0] regs_8_io_in;
  wire [63:0] regs_8_io_init;
  wire [63:0] regs_8_io_out;
  wire  regs_8_io_enable;
  wire  regs_9_clock;
  wire  regs_9_reset;
  wire [63:0] regs_9_io_in;
  wire [63:0] regs_9_io_init;
  wire [63:0] regs_9_io_out;
  wire  regs_9_io_enable;
  wire  regs_10_clock;
  wire  regs_10_reset;
  wire [63:0] regs_10_io_in;
  wire [63:0] regs_10_io_init;
  wire [63:0] regs_10_io_out;
  wire  regs_10_io_enable;
  wire  regs_11_clock;
  wire  regs_11_reset;
  wire [63:0] regs_11_io_in;
  wire [63:0] regs_11_io_init;
  wire [63:0] regs_11_io_out;
  wire  regs_11_io_enable;
  wire  regs_12_clock;
  wire  regs_12_reset;
  wire [63:0] regs_12_io_in;
  wire [63:0] regs_12_io_init;
  wire [63:0] regs_12_io_out;
  wire  regs_12_io_enable;
  wire  regs_13_clock;
  wire  regs_13_reset;
  wire [63:0] regs_13_io_in;
  wire [63:0] regs_13_io_init;
  wire [63:0] regs_13_io_out;
  wire  regs_13_io_enable;
  wire  regs_14_clock;
  wire  regs_14_reset;
  wire [63:0] regs_14_io_in;
  wire [63:0] regs_14_io_init;
  wire [63:0] regs_14_io_out;
  wire  regs_14_io_enable;
  wire  regs_15_clock;
  wire  regs_15_reset;
  wire [63:0] regs_15_io_in;
  wire [63:0] regs_15_io_init;
  wire [63:0] regs_15_io_out;
  wire  regs_15_io_enable;
  wire  regs_16_clock;
  wire  regs_16_reset;
  wire [63:0] regs_16_io_in;
  wire [63:0] regs_16_io_init;
  wire [63:0] regs_16_io_out;
  wire  regs_16_io_enable;
  wire  regs_17_clock;
  wire  regs_17_reset;
  wire [63:0] regs_17_io_in;
  wire [63:0] regs_17_io_init;
  wire [63:0] regs_17_io_out;
  wire  regs_17_io_enable;
  wire  regs_18_clock;
  wire  regs_18_reset;
  wire [63:0] regs_18_io_in;
  wire [63:0] regs_18_io_init;
  wire [63:0] regs_18_io_out;
  wire  regs_18_io_enable;
  wire  regs_19_clock;
  wire  regs_19_reset;
  wire [63:0] regs_19_io_in;
  wire [63:0] regs_19_io_init;
  wire [63:0] regs_19_io_out;
  wire  regs_19_io_enable;
  wire  regs_20_clock;
  wire  regs_20_reset;
  wire [63:0] regs_20_io_in;
  wire [63:0] regs_20_io_init;
  wire [63:0] regs_20_io_out;
  wire  regs_20_io_enable;
  wire  regs_21_clock;
  wire  regs_21_reset;
  wire [63:0] regs_21_io_in;
  wire [63:0] regs_21_io_init;
  wire [63:0] regs_21_io_out;
  wire  regs_21_io_enable;
  wire  regs_22_clock;
  wire  regs_22_reset;
  wire [63:0] regs_22_io_in;
  wire [63:0] regs_22_io_init;
  wire [63:0] regs_22_io_out;
  wire  regs_22_io_enable;
  wire  regs_23_clock;
  wire  regs_23_reset;
  wire [63:0] regs_23_io_in;
  wire [63:0] regs_23_io_init;
  wire [63:0] regs_23_io_out;
  wire  regs_23_io_enable;
  wire  regs_24_clock;
  wire  regs_24_reset;
  wire [63:0] regs_24_io_in;
  wire [63:0] regs_24_io_init;
  wire [63:0] regs_24_io_out;
  wire  regs_24_io_enable;
  wire  regs_25_clock;
  wire  regs_25_reset;
  wire [63:0] regs_25_io_in;
  wire [63:0] regs_25_io_init;
  wire [63:0] regs_25_io_out;
  wire  regs_25_io_enable;
  wire  regs_26_clock;
  wire  regs_26_reset;
  wire [63:0] regs_26_io_in;
  wire [63:0] regs_26_io_init;
  wire [63:0] regs_26_io_out;
  wire  regs_26_io_enable;
  wire  regs_27_clock;
  wire  regs_27_reset;
  wire [63:0] regs_27_io_in;
  wire [63:0] regs_27_io_init;
  wire [63:0] regs_27_io_out;
  wire  regs_27_io_enable;
  wire  regs_28_clock;
  wire  regs_28_reset;
  wire [63:0] regs_28_io_in;
  wire [63:0] regs_28_io_init;
  wire [63:0] regs_28_io_out;
  wire  regs_28_io_enable;
  wire  regs_29_clock;
  wire  regs_29_reset;
  wire [63:0] regs_29_io_in;
  wire [63:0] regs_29_io_init;
  wire [63:0] regs_29_io_out;
  wire  regs_29_io_enable;
  wire  regs_30_clock;
  wire  regs_30_reset;
  wire [63:0] regs_30_io_in;
  wire [63:0] regs_30_io_init;
  wire [63:0] regs_30_io_out;
  wire  regs_30_io_enable;
  wire  regs_31_clock;
  wire  regs_31_reset;
  wire [63:0] regs_31_io_in;
  wire [63:0] regs_31_io_init;
  wire [63:0] regs_31_io_out;
  wire  regs_31_io_enable;
  wire  regs_32_clock;
  wire  regs_32_reset;
  wire [63:0] regs_32_io_in;
  wire [63:0] regs_32_io_init;
  wire [63:0] regs_32_io_out;
  wire  regs_32_io_enable;
  wire  regs_33_clock;
  wire  regs_33_reset;
  wire [63:0] regs_33_io_in;
  wire [63:0] regs_33_io_init;
  wire [63:0] regs_33_io_out;
  wire  regs_33_io_enable;
  wire  regs_34_clock;
  wire  regs_34_reset;
  wire [63:0] regs_34_io_in;
  wire [63:0] regs_34_io_init;
  wire [63:0] regs_34_io_out;
  wire  regs_34_io_enable;
  wire  regs_35_clock;
  wire  regs_35_reset;
  wire [63:0] regs_35_io_in;
  wire [63:0] regs_35_io_init;
  wire [63:0] regs_35_io_out;
  wire  regs_35_io_enable;
  wire  regs_36_clock;
  wire  regs_36_reset;
  wire [63:0] regs_36_io_in;
  wire [63:0] regs_36_io_init;
  wire [63:0] regs_36_io_out;
  wire  regs_36_io_enable;
  wire  regs_37_clock;
  wire  regs_37_reset;
  wire [63:0] regs_37_io_in;
  wire [63:0] regs_37_io_init;
  wire [63:0] regs_37_io_out;
  wire  regs_37_io_enable;
  wire  regs_38_clock;
  wire  regs_38_reset;
  wire [63:0] regs_38_io_in;
  wire [63:0] regs_38_io_init;
  wire [63:0] regs_38_io_out;
  wire  regs_38_io_enable;
  wire  regs_39_clock;
  wire  regs_39_reset;
  wire [63:0] regs_39_io_in;
  wire [63:0] regs_39_io_init;
  wire [63:0] regs_39_io_out;
  wire  regs_39_io_enable;
  wire  regs_40_clock;
  wire  regs_40_reset;
  wire [63:0] regs_40_io_in;
  wire [63:0] regs_40_io_init;
  wire [63:0] regs_40_io_out;
  wire  regs_40_io_enable;
  wire  regs_41_clock;
  wire  regs_41_reset;
  wire [63:0] regs_41_io_in;
  wire [63:0] regs_41_io_init;
  wire [63:0] regs_41_io_out;
  wire  regs_41_io_enable;
  wire  regs_42_clock;
  wire  regs_42_reset;
  wire [63:0] regs_42_io_in;
  wire [63:0] regs_42_io_init;
  wire [63:0] regs_42_io_out;
  wire  regs_42_io_enable;
  wire  regs_43_clock;
  wire  regs_43_reset;
  wire [63:0] regs_43_io_in;
  wire [63:0] regs_43_io_init;
  wire [63:0] regs_43_io_out;
  wire  regs_43_io_enable;
  wire  regs_44_clock;
  wire  regs_44_reset;
  wire [63:0] regs_44_io_in;
  wire [63:0] regs_44_io_init;
  wire [63:0] regs_44_io_out;
  wire  regs_44_io_enable;
  wire  regs_45_clock;
  wire  regs_45_reset;
  wire [63:0] regs_45_io_in;
  wire [63:0] regs_45_io_init;
  wire [63:0] regs_45_io_out;
  wire  regs_45_io_enable;
  wire  regs_46_clock;
  wire  regs_46_reset;
  wire [63:0] regs_46_io_in;
  wire [63:0] regs_46_io_init;
  wire [63:0] regs_46_io_out;
  wire  regs_46_io_enable;
  wire  regs_47_clock;
  wire  regs_47_reset;
  wire [63:0] regs_47_io_in;
  wire [63:0] regs_47_io_init;
  wire [63:0] regs_47_io_out;
  wire  regs_47_io_enable;
  wire  regs_48_clock;
  wire  regs_48_reset;
  wire [63:0] regs_48_io_in;
  wire [63:0] regs_48_io_init;
  wire [63:0] regs_48_io_out;
  wire  regs_48_io_enable;
  wire  regs_49_clock;
  wire  regs_49_reset;
  wire [63:0] regs_49_io_in;
  wire [63:0] regs_49_io_init;
  wire [63:0] regs_49_io_out;
  wire  regs_49_io_enable;
  wire  regs_50_clock;
  wire  regs_50_reset;
  wire [63:0] regs_50_io_in;
  wire [63:0] regs_50_io_init;
  wire [63:0] regs_50_io_out;
  wire  regs_50_io_enable;
  wire  regs_51_clock;
  wire  regs_51_reset;
  wire [63:0] regs_51_io_in;
  wire [63:0] regs_51_io_init;
  wire [63:0] regs_51_io_out;
  wire  regs_51_io_enable;
  wire  regs_52_clock;
  wire  regs_52_reset;
  wire [63:0] regs_52_io_in;
  wire [63:0] regs_52_io_init;
  wire [63:0] regs_52_io_out;
  wire  regs_52_io_enable;
  wire  regs_53_clock;
  wire  regs_53_reset;
  wire [63:0] regs_53_io_in;
  wire [63:0] regs_53_io_init;
  wire [63:0] regs_53_io_out;
  wire  regs_53_io_enable;
  wire  regs_54_clock;
  wire  regs_54_reset;
  wire [63:0] regs_54_io_in;
  wire [63:0] regs_54_io_init;
  wire [63:0] regs_54_io_out;
  wire  regs_54_io_enable;
  wire  regs_55_clock;
  wire  regs_55_reset;
  wire [63:0] regs_55_io_in;
  wire [63:0] regs_55_io_init;
  wire [63:0] regs_55_io_out;
  wire  regs_55_io_enable;
  wire  regs_56_clock;
  wire  regs_56_reset;
  wire [63:0] regs_56_io_in;
  wire [63:0] regs_56_io_init;
  wire [63:0] regs_56_io_out;
  wire  regs_56_io_enable;
  wire  regs_57_clock;
  wire  regs_57_reset;
  wire [63:0] regs_57_io_in;
  wire [63:0] regs_57_io_init;
  wire [63:0] regs_57_io_out;
  wire  regs_57_io_enable;
  wire  regs_58_clock;
  wire  regs_58_reset;
  wire [63:0] regs_58_io_in;
  wire [63:0] regs_58_io_init;
  wire [63:0] regs_58_io_out;
  wire  regs_58_io_enable;
  wire  regs_59_clock;
  wire  regs_59_reset;
  wire [63:0] regs_59_io_in;
  wire [63:0] regs_59_io_init;
  wire [63:0] regs_59_io_out;
  wire  regs_59_io_enable;
  wire  regs_60_clock;
  wire  regs_60_reset;
  wire [63:0] regs_60_io_in;
  wire [63:0] regs_60_io_init;
  wire [63:0] regs_60_io_out;
  wire  regs_60_io_enable;
  wire  regs_61_clock;
  wire  regs_61_reset;
  wire [63:0] regs_61_io_in;
  wire [63:0] regs_61_io_init;
  wire [63:0] regs_61_io_out;
  wire  regs_61_io_enable;
  wire  regs_62_clock;
  wire  regs_62_reset;
  wire [63:0] regs_62_io_in;
  wire [63:0] regs_62_io_init;
  wire [63:0] regs_62_io_out;
  wire  regs_62_io_enable;
  wire  regs_63_clock;
  wire  regs_63_reset;
  wire [63:0] regs_63_io_in;
  wire [63:0] regs_63_io_init;
  wire [63:0] regs_63_io_out;
  wire  regs_63_io_enable;
  wire  regs_64_clock;
  wire  regs_64_reset;
  wire [63:0] regs_64_io_in;
  wire [63:0] regs_64_io_init;
  wire [63:0] regs_64_io_out;
  wire  regs_64_io_enable;
  wire  regs_65_clock;
  wire  regs_65_reset;
  wire [63:0] regs_65_io_in;
  wire [63:0] regs_65_io_init;
  wire [63:0] regs_65_io_out;
  wire  regs_65_io_enable;
  wire  regs_66_clock;
  wire  regs_66_reset;
  wire [63:0] regs_66_io_in;
  wire [63:0] regs_66_io_init;
  wire [63:0] regs_66_io_out;
  wire  regs_66_io_enable;
  wire  regs_67_clock;
  wire  regs_67_reset;
  wire [63:0] regs_67_io_in;
  wire [63:0] regs_67_io_init;
  wire [63:0] regs_67_io_out;
  wire  regs_67_io_enable;
  wire  regs_68_clock;
  wire  regs_68_reset;
  wire [63:0] regs_68_io_in;
  wire [63:0] regs_68_io_init;
  wire [63:0] regs_68_io_out;
  wire  regs_68_io_enable;
  wire  regs_69_clock;
  wire  regs_69_reset;
  wire [63:0] regs_69_io_in;
  wire [63:0] regs_69_io_init;
  wire [63:0] regs_69_io_out;
  wire  regs_69_io_enable;
  wire  regs_70_clock;
  wire  regs_70_reset;
  wire [63:0] regs_70_io_in;
  wire [63:0] regs_70_io_init;
  wire [63:0] regs_70_io_out;
  wire  regs_70_io_enable;
  wire  regs_71_clock;
  wire  regs_71_reset;
  wire [63:0] regs_71_io_in;
  wire [63:0] regs_71_io_init;
  wire [63:0] regs_71_io_out;
  wire  regs_71_io_enable;
  wire  regs_72_clock;
  wire  regs_72_reset;
  wire [63:0] regs_72_io_in;
  wire [63:0] regs_72_io_init;
  wire [63:0] regs_72_io_out;
  wire  regs_72_io_enable;
  wire  regs_73_clock;
  wire  regs_73_reset;
  wire [63:0] regs_73_io_in;
  wire [63:0] regs_73_io_init;
  wire [63:0] regs_73_io_out;
  wire  regs_73_io_enable;
  wire  regs_74_clock;
  wire  regs_74_reset;
  wire [63:0] regs_74_io_in;
  wire [63:0] regs_74_io_init;
  wire [63:0] regs_74_io_out;
  wire  regs_74_io_enable;
  wire  regs_75_clock;
  wire  regs_75_reset;
  wire [63:0] regs_75_io_in;
  wire [63:0] regs_75_io_init;
  wire [63:0] regs_75_io_out;
  wire  regs_75_io_enable;
  wire  regs_76_clock;
  wire  regs_76_reset;
  wire [63:0] regs_76_io_in;
  wire [63:0] regs_76_io_init;
  wire [63:0] regs_76_io_out;
  wire  regs_76_io_enable;
  wire  regs_77_clock;
  wire  regs_77_reset;
  wire [63:0] regs_77_io_in;
  wire [63:0] regs_77_io_init;
  wire [63:0] regs_77_io_out;
  wire  regs_77_io_enable;
  wire  regs_78_clock;
  wire  regs_78_reset;
  wire [63:0] regs_78_io_in;
  wire [63:0] regs_78_io_init;
  wire [63:0] regs_78_io_out;
  wire  regs_78_io_enable;
  wire  regs_79_clock;
  wire  regs_79_reset;
  wire [63:0] regs_79_io_in;
  wire [63:0] regs_79_io_init;
  wire [63:0] regs_79_io_out;
  wire  regs_79_io_enable;
  wire  regs_80_clock;
  wire  regs_80_reset;
  wire [63:0] regs_80_io_in;
  wire [63:0] regs_80_io_init;
  wire [63:0] regs_80_io_out;
  wire  regs_80_io_enable;
  wire  regs_81_clock;
  wire  regs_81_reset;
  wire [63:0] regs_81_io_in;
  wire [63:0] regs_81_io_init;
  wire [63:0] regs_81_io_out;
  wire  regs_81_io_enable;
  wire  regs_82_clock;
  wire  regs_82_reset;
  wire [63:0] regs_82_io_in;
  wire [63:0] regs_82_io_init;
  wire [63:0] regs_82_io_out;
  wire  regs_82_io_enable;
  wire  regs_83_clock;
  wire  regs_83_reset;
  wire [63:0] regs_83_io_in;
  wire [63:0] regs_83_io_init;
  wire [63:0] regs_83_io_out;
  wire  regs_83_io_enable;
  wire  regs_84_clock;
  wire  regs_84_reset;
  wire [63:0] regs_84_io_in;
  wire [63:0] regs_84_io_init;
  wire [63:0] regs_84_io_out;
  wire  regs_84_io_enable;
  wire  regs_85_clock;
  wire  regs_85_reset;
  wire [63:0] regs_85_io_in;
  wire [63:0] regs_85_io_init;
  wire [63:0] regs_85_io_out;
  wire  regs_85_io_enable;
  wire  regs_86_clock;
  wire  regs_86_reset;
  wire [63:0] regs_86_io_in;
  wire [63:0] regs_86_io_init;
  wire [63:0] regs_86_io_out;
  wire  regs_86_io_enable;
  wire  regs_87_clock;
  wire  regs_87_reset;
  wire [63:0] regs_87_io_in;
  wire [63:0] regs_87_io_init;
  wire [63:0] regs_87_io_out;
  wire  regs_87_io_enable;
  wire  regs_88_clock;
  wire  regs_88_reset;
  wire [63:0] regs_88_io_in;
  wire [63:0] regs_88_io_init;
  wire [63:0] regs_88_io_out;
  wire  regs_88_io_enable;
  wire  regs_89_clock;
  wire  regs_89_reset;
  wire [63:0] regs_89_io_in;
  wire [63:0] regs_89_io_init;
  wire [63:0] regs_89_io_out;
  wire  regs_89_io_enable;
  wire  regs_90_clock;
  wire  regs_90_reset;
  wire [63:0] regs_90_io_in;
  wire [63:0] regs_90_io_init;
  wire [63:0] regs_90_io_out;
  wire  regs_90_io_enable;
  wire  regs_91_clock;
  wire  regs_91_reset;
  wire [63:0] regs_91_io_in;
  wire [63:0] regs_91_io_init;
  wire [63:0] regs_91_io_out;
  wire  regs_91_io_enable;
  wire  regs_92_clock;
  wire  regs_92_reset;
  wire [63:0] regs_92_io_in;
  wire [63:0] regs_92_io_init;
  wire [63:0] regs_92_io_out;
  wire  regs_92_io_enable;
  wire  regs_93_clock;
  wire  regs_93_reset;
  wire [63:0] regs_93_io_in;
  wire [63:0] regs_93_io_init;
  wire [63:0] regs_93_io_out;
  wire  regs_93_io_enable;
  wire  regs_94_clock;
  wire  regs_94_reset;
  wire [63:0] regs_94_io_in;
  wire [63:0] regs_94_io_init;
  wire [63:0] regs_94_io_out;
  wire  regs_94_io_enable;
  wire  regs_95_clock;
  wire  regs_95_reset;
  wire [63:0] regs_95_io_in;
  wire [63:0] regs_95_io_init;
  wire [63:0] regs_95_io_out;
  wire  regs_95_io_enable;
  wire  regs_96_clock;
  wire  regs_96_reset;
  wire [63:0] regs_96_io_in;
  wire [63:0] regs_96_io_init;
  wire [63:0] regs_96_io_out;
  wire  regs_96_io_enable;
  wire  regs_97_clock;
  wire  regs_97_reset;
  wire [63:0] regs_97_io_in;
  wire [63:0] regs_97_io_init;
  wire [63:0] regs_97_io_out;
  wire  regs_97_io_enable;
  wire  regs_98_clock;
  wire  regs_98_reset;
  wire [63:0] regs_98_io_in;
  wire [63:0] regs_98_io_init;
  wire [63:0] regs_98_io_out;
  wire  regs_98_io_enable;
  wire  regs_99_clock;
  wire  regs_99_reset;
  wire [63:0] regs_99_io_in;
  wire [63:0] regs_99_io_init;
  wire [63:0] regs_99_io_out;
  wire  regs_99_io_enable;
  wire  regs_100_clock;
  wire  regs_100_reset;
  wire [63:0] regs_100_io_in;
  wire [63:0] regs_100_io_init;
  wire [63:0] regs_100_io_out;
  wire  regs_100_io_enable;
  wire  regs_101_clock;
  wire  regs_101_reset;
  wire [63:0] regs_101_io_in;
  wire [63:0] regs_101_io_init;
  wire [63:0] regs_101_io_out;
  wire  regs_101_io_enable;
  wire  regs_102_clock;
  wire  regs_102_reset;
  wire [63:0] regs_102_io_in;
  wire [63:0] regs_102_io_init;
  wire [63:0] regs_102_io_out;
  wire  regs_102_io_enable;
  wire  regs_103_clock;
  wire  regs_103_reset;
  wire [63:0] regs_103_io_in;
  wire [63:0] regs_103_io_init;
  wire [63:0] regs_103_io_out;
  wire  regs_103_io_enable;
  wire  regs_104_clock;
  wire  regs_104_reset;
  wire [63:0] regs_104_io_in;
  wire [63:0] regs_104_io_init;
  wire [63:0] regs_104_io_out;
  wire  regs_104_io_enable;
  wire  regs_105_clock;
  wire  regs_105_reset;
  wire [63:0] regs_105_io_in;
  wire [63:0] regs_105_io_init;
  wire [63:0] regs_105_io_out;
  wire  regs_105_io_enable;
  wire  regs_106_clock;
  wire  regs_106_reset;
  wire [63:0] regs_106_io_in;
  wire [63:0] regs_106_io_init;
  wire [63:0] regs_106_io_out;
  wire  regs_106_io_enable;
  wire  regs_107_clock;
  wire  regs_107_reset;
  wire [63:0] regs_107_io_in;
  wire [63:0] regs_107_io_init;
  wire [63:0] regs_107_io_out;
  wire  regs_107_io_enable;
  wire  regs_108_clock;
  wire  regs_108_reset;
  wire [63:0] regs_108_io_in;
  wire [63:0] regs_108_io_init;
  wire [63:0] regs_108_io_out;
  wire  regs_108_io_enable;
  wire  regs_109_clock;
  wire  regs_109_reset;
  wire [63:0] regs_109_io_in;
  wire [63:0] regs_109_io_init;
  wire [63:0] regs_109_io_out;
  wire  regs_109_io_enable;
  wire  regs_110_clock;
  wire  regs_110_reset;
  wire [63:0] regs_110_io_in;
  wire [63:0] regs_110_io_init;
  wire [63:0] regs_110_io_out;
  wire  regs_110_io_enable;
  wire  regs_111_clock;
  wire  regs_111_reset;
  wire [63:0] regs_111_io_in;
  wire [63:0] regs_111_io_init;
  wire [63:0] regs_111_io_out;
  wire  regs_111_io_enable;
  wire  regs_112_clock;
  wire  regs_112_reset;
  wire [63:0] regs_112_io_in;
  wire [63:0] regs_112_io_init;
  wire [63:0] regs_112_io_out;
  wire  regs_112_io_enable;
  wire  regs_113_clock;
  wire  regs_113_reset;
  wire [63:0] regs_113_io_in;
  wire [63:0] regs_113_io_init;
  wire [63:0] regs_113_io_out;
  wire  regs_113_io_enable;
  wire  regs_114_clock;
  wire  regs_114_reset;
  wire [63:0] regs_114_io_in;
  wire [63:0] regs_114_io_init;
  wire [63:0] regs_114_io_out;
  wire  regs_114_io_enable;
  wire  regs_115_clock;
  wire  regs_115_reset;
  wire [63:0] regs_115_io_in;
  wire [63:0] regs_115_io_init;
  wire [63:0] regs_115_io_out;
  wire  regs_115_io_enable;
  wire  regs_116_clock;
  wire  regs_116_reset;
  wire [63:0] regs_116_io_in;
  wire [63:0] regs_116_io_init;
  wire [63:0] regs_116_io_out;
  wire  regs_116_io_enable;
  wire  regs_117_clock;
  wire  regs_117_reset;
  wire [63:0] regs_117_io_in;
  wire [63:0] regs_117_io_init;
  wire [63:0] regs_117_io_out;
  wire  regs_117_io_enable;
  wire  regs_118_clock;
  wire  regs_118_reset;
  wire [63:0] regs_118_io_in;
  wire [63:0] regs_118_io_init;
  wire [63:0] regs_118_io_out;
  wire  regs_118_io_enable;
  wire  regs_119_clock;
  wire  regs_119_reset;
  wire [63:0] regs_119_io_in;
  wire [63:0] regs_119_io_init;
  wire [63:0] regs_119_io_out;
  wire  regs_119_io_enable;
  wire  regs_120_clock;
  wire  regs_120_reset;
  wire [63:0] regs_120_io_in;
  wire [63:0] regs_120_io_init;
  wire [63:0] regs_120_io_out;
  wire  regs_120_io_enable;
  wire  regs_121_clock;
  wire  regs_121_reset;
  wire [63:0] regs_121_io_in;
  wire [63:0] regs_121_io_init;
  wire [63:0] regs_121_io_out;
  wire  regs_121_io_enable;
  wire  regs_122_clock;
  wire  regs_122_reset;
  wire [63:0] regs_122_io_in;
  wire [63:0] regs_122_io_init;
  wire [63:0] regs_122_io_out;
  wire  regs_122_io_enable;
  wire  regs_123_clock;
  wire  regs_123_reset;
  wire [63:0] regs_123_io_in;
  wire [63:0] regs_123_io_init;
  wire [63:0] regs_123_io_out;
  wire  regs_123_io_enable;
  wire  regs_124_clock;
  wire  regs_124_reset;
  wire [63:0] regs_124_io_in;
  wire [63:0] regs_124_io_init;
  wire [63:0] regs_124_io_out;
  wire  regs_124_io_enable;
  wire  regs_125_clock;
  wire  regs_125_reset;
  wire [63:0] regs_125_io_in;
  wire [63:0] regs_125_io_init;
  wire [63:0] regs_125_io_out;
  wire  regs_125_io_enable;
  wire  regs_126_clock;
  wire  regs_126_reset;
  wire [63:0] regs_126_io_in;
  wire [63:0] regs_126_io_init;
  wire [63:0] regs_126_io_out;
  wire  regs_126_io_enable;
  wire  regs_127_clock;
  wire  regs_127_reset;
  wire [63:0] regs_127_io_in;
  wire [63:0] regs_127_io_init;
  wire [63:0] regs_127_io_out;
  wire  regs_127_io_enable;
  wire  regs_128_clock;
  wire  regs_128_reset;
  wire [63:0] regs_128_io_in;
  wire [63:0] regs_128_io_init;
  wire [63:0] regs_128_io_out;
  wire  regs_128_io_enable;
  wire  regs_129_clock;
  wire  regs_129_reset;
  wire [63:0] regs_129_io_in;
  wire [63:0] regs_129_io_init;
  wire [63:0] regs_129_io_out;
  wire  regs_129_io_enable;
  wire  regs_130_clock;
  wire  regs_130_reset;
  wire [63:0] regs_130_io_in;
  wire [63:0] regs_130_io_init;
  wire [63:0] regs_130_io_out;
  wire  regs_130_io_enable;
  wire  regs_131_clock;
  wire  regs_131_reset;
  wire [63:0] regs_131_io_in;
  wire [63:0] regs_131_io_init;
  wire [63:0] regs_131_io_out;
  wire  regs_131_io_enable;
  wire  regs_132_clock;
  wire  regs_132_reset;
  wire [63:0] regs_132_io_in;
  wire [63:0] regs_132_io_init;
  wire [63:0] regs_132_io_out;
  wire  regs_132_io_enable;
  wire  regs_133_clock;
  wire  regs_133_reset;
  wire [63:0] regs_133_io_in;
  wire [63:0] regs_133_io_init;
  wire [63:0] regs_133_io_out;
  wire  regs_133_io_enable;
  wire  regs_134_clock;
  wire  regs_134_reset;
  wire [63:0] regs_134_io_in;
  wire [63:0] regs_134_io_init;
  wire [63:0] regs_134_io_out;
  wire  regs_134_io_enable;
  wire  regs_135_clock;
  wire  regs_135_reset;
  wire [63:0] regs_135_io_in;
  wire [63:0] regs_135_io_init;
  wire [63:0] regs_135_io_out;
  wire  regs_135_io_enable;
  wire  regs_136_clock;
  wire  regs_136_reset;
  wire [63:0] regs_136_io_in;
  wire [63:0] regs_136_io_init;
  wire [63:0] regs_136_io_out;
  wire  regs_136_io_enable;
  wire  regs_137_clock;
  wire  regs_137_reset;
  wire [63:0] regs_137_io_in;
  wire [63:0] regs_137_io_init;
  wire [63:0] regs_137_io_out;
  wire  regs_137_io_enable;
  wire  regs_138_clock;
  wire  regs_138_reset;
  wire [63:0] regs_138_io_in;
  wire [63:0] regs_138_io_init;
  wire [63:0] regs_138_io_out;
  wire  regs_138_io_enable;
  wire  regs_139_clock;
  wire  regs_139_reset;
  wire [63:0] regs_139_io_in;
  wire [63:0] regs_139_io_init;
  wire [63:0] regs_139_io_out;
  wire  regs_139_io_enable;
  wire  regs_140_clock;
  wire  regs_140_reset;
  wire [63:0] regs_140_io_in;
  wire [63:0] regs_140_io_init;
  wire [63:0] regs_140_io_out;
  wire  regs_140_io_enable;
  wire  regs_141_clock;
  wire  regs_141_reset;
  wire [63:0] regs_141_io_in;
  wire [63:0] regs_141_io_init;
  wire [63:0] regs_141_io_out;
  wire  regs_141_io_enable;
  wire  regs_142_clock;
  wire  regs_142_reset;
  wire [63:0] regs_142_io_in;
  wire [63:0] regs_142_io_init;
  wire [63:0] regs_142_io_out;
  wire  regs_142_io_enable;
  wire  regs_143_clock;
  wire  regs_143_reset;
  wire [63:0] regs_143_io_in;
  wire [63:0] regs_143_io_init;
  wire [63:0] regs_143_io_out;
  wire  regs_143_io_enable;
  wire  regs_144_clock;
  wire  regs_144_reset;
  wire [63:0] regs_144_io_in;
  wire [63:0] regs_144_io_init;
  wire [63:0] regs_144_io_out;
  wire  regs_144_io_enable;
  wire  regs_145_clock;
  wire  regs_145_reset;
  wire [63:0] regs_145_io_in;
  wire [63:0] regs_145_io_init;
  wire [63:0] regs_145_io_out;
  wire  regs_145_io_enable;
  wire  regs_146_clock;
  wire  regs_146_reset;
  wire [63:0] regs_146_io_in;
  wire [63:0] regs_146_io_init;
  wire [63:0] regs_146_io_out;
  wire  regs_146_io_enable;
  wire  regs_147_clock;
  wire  regs_147_reset;
  wire [63:0] regs_147_io_in;
  wire [63:0] regs_147_io_init;
  wire [63:0] regs_147_io_out;
  wire  regs_147_io_enable;
  wire  regs_148_clock;
  wire  regs_148_reset;
  wire [63:0] regs_148_io_in;
  wire [63:0] regs_148_io_init;
  wire [63:0] regs_148_io_out;
  wire  regs_148_io_enable;
  wire  regs_149_clock;
  wire  regs_149_reset;
  wire [63:0] regs_149_io_in;
  wire [63:0] regs_149_io_init;
  wire [63:0] regs_149_io_out;
  wire  regs_149_io_enable;
  wire  regs_150_clock;
  wire  regs_150_reset;
  wire [63:0] regs_150_io_in;
  wire [63:0] regs_150_io_init;
  wire [63:0] regs_150_io_out;
  wire  regs_150_io_enable;
  wire  regs_151_clock;
  wire  regs_151_reset;
  wire [63:0] regs_151_io_in;
  wire [63:0] regs_151_io_init;
  wire [63:0] regs_151_io_out;
  wire  regs_151_io_enable;
  wire  regs_152_clock;
  wire  regs_152_reset;
  wire [63:0] regs_152_io_in;
  wire [63:0] regs_152_io_init;
  wire [63:0] regs_152_io_out;
  wire  regs_152_io_enable;
  wire  regs_153_clock;
  wire  regs_153_reset;
  wire [63:0] regs_153_io_in;
  wire [63:0] regs_153_io_init;
  wire [63:0] regs_153_io_out;
  wire  regs_153_io_enable;
  wire  regs_154_clock;
  wire  regs_154_reset;
  wire [63:0] regs_154_io_in;
  wire [63:0] regs_154_io_init;
  wire [63:0] regs_154_io_out;
  wire  regs_154_io_enable;
  wire  regs_155_clock;
  wire  regs_155_reset;
  wire [63:0] regs_155_io_in;
  wire [63:0] regs_155_io_init;
  wire [63:0] regs_155_io_out;
  wire  regs_155_io_enable;
  wire  regs_156_clock;
  wire  regs_156_reset;
  wire [63:0] regs_156_io_in;
  wire [63:0] regs_156_io_init;
  wire [63:0] regs_156_io_out;
  wire  regs_156_io_enable;
  wire  regs_157_clock;
  wire  regs_157_reset;
  wire [63:0] regs_157_io_in;
  wire [63:0] regs_157_io_init;
  wire [63:0] regs_157_io_out;
  wire  regs_157_io_enable;
  wire  regs_158_clock;
  wire  regs_158_reset;
  wire [63:0] regs_158_io_in;
  wire [63:0] regs_158_io_init;
  wire [63:0] regs_158_io_out;
  wire  regs_158_io_enable;
  wire  regs_159_clock;
  wire  regs_159_reset;
  wire [63:0] regs_159_io_in;
  wire [63:0] regs_159_io_init;
  wire [63:0] regs_159_io_out;
  wire  regs_159_io_enable;
  wire  regs_160_clock;
  wire  regs_160_reset;
  wire [63:0] regs_160_io_in;
  wire [63:0] regs_160_io_init;
  wire [63:0] regs_160_io_out;
  wire  regs_160_io_enable;
  wire  regs_161_clock;
  wire  regs_161_reset;
  wire [63:0] regs_161_io_in;
  wire [63:0] regs_161_io_init;
  wire [63:0] regs_161_io_out;
  wire  regs_161_io_enable;
  wire  regs_162_clock;
  wire  regs_162_reset;
  wire [63:0] regs_162_io_in;
  wire [63:0] regs_162_io_init;
  wire [63:0] regs_162_io_out;
  wire  regs_162_io_enable;
  wire  regs_163_clock;
  wire  regs_163_reset;
  wire [63:0] regs_163_io_in;
  wire [63:0] regs_163_io_init;
  wire [63:0] regs_163_io_out;
  wire  regs_163_io_enable;
  wire  regs_164_clock;
  wire  regs_164_reset;
  wire [63:0] regs_164_io_in;
  wire [63:0] regs_164_io_init;
  wire [63:0] regs_164_io_out;
  wire  regs_164_io_enable;
  wire  regs_165_clock;
  wire  regs_165_reset;
  wire [63:0] regs_165_io_in;
  wire [63:0] regs_165_io_init;
  wire [63:0] regs_165_io_out;
  wire  regs_165_io_enable;
  wire  regs_166_clock;
  wire  regs_166_reset;
  wire [63:0] regs_166_io_in;
  wire [63:0] regs_166_io_init;
  wire [63:0] regs_166_io_out;
  wire  regs_166_io_enable;
  wire  regs_167_clock;
  wire  regs_167_reset;
  wire [63:0] regs_167_io_in;
  wire [63:0] regs_167_io_init;
  wire [63:0] regs_167_io_out;
  wire  regs_167_io_enable;
  wire  regs_168_clock;
  wire  regs_168_reset;
  wire [63:0] regs_168_io_in;
  wire [63:0] regs_168_io_init;
  wire [63:0] regs_168_io_out;
  wire  regs_168_io_enable;
  wire  regs_169_clock;
  wire  regs_169_reset;
  wire [63:0] regs_169_io_in;
  wire [63:0] regs_169_io_init;
  wire [63:0] regs_169_io_out;
  wire  regs_169_io_enable;
  wire  regs_170_clock;
  wire  regs_170_reset;
  wire [63:0] regs_170_io_in;
  wire [63:0] regs_170_io_init;
  wire [63:0] regs_170_io_out;
  wire  regs_170_io_enable;
  wire  regs_171_clock;
  wire  regs_171_reset;
  wire [63:0] regs_171_io_in;
  wire [63:0] regs_171_io_init;
  wire [63:0] regs_171_io_out;
  wire  regs_171_io_enable;
  wire  regs_172_clock;
  wire  regs_172_reset;
  wire [63:0] regs_172_io_in;
  wire [63:0] regs_172_io_init;
  wire [63:0] regs_172_io_out;
  wire  regs_172_io_enable;
  wire  regs_173_clock;
  wire  regs_173_reset;
  wire [63:0] regs_173_io_in;
  wire [63:0] regs_173_io_init;
  wire [63:0] regs_173_io_out;
  wire  regs_173_io_enable;
  wire  regs_174_clock;
  wire  regs_174_reset;
  wire [63:0] regs_174_io_in;
  wire [63:0] regs_174_io_init;
  wire [63:0] regs_174_io_out;
  wire  regs_174_io_enable;
  wire  regs_175_clock;
  wire  regs_175_reset;
  wire [63:0] regs_175_io_in;
  wire [63:0] regs_175_io_init;
  wire [63:0] regs_175_io_out;
  wire  regs_175_io_enable;
  wire  regs_176_clock;
  wire  regs_176_reset;
  wire [63:0] regs_176_io_in;
  wire [63:0] regs_176_io_init;
  wire [63:0] regs_176_io_out;
  wire  regs_176_io_enable;
  wire  regs_177_clock;
  wire  regs_177_reset;
  wire [63:0] regs_177_io_in;
  wire [63:0] regs_177_io_init;
  wire [63:0] regs_177_io_out;
  wire  regs_177_io_enable;
  wire  regs_178_clock;
  wire  regs_178_reset;
  wire [63:0] regs_178_io_in;
  wire [63:0] regs_178_io_init;
  wire [63:0] regs_178_io_out;
  wire  regs_178_io_enable;
  wire  regs_179_clock;
  wire  regs_179_reset;
  wire [63:0] regs_179_io_in;
  wire [63:0] regs_179_io_init;
  wire [63:0] regs_179_io_out;
  wire  regs_179_io_enable;
  wire  regs_180_clock;
  wire  regs_180_reset;
  wire [63:0] regs_180_io_in;
  wire [63:0] regs_180_io_init;
  wire [63:0] regs_180_io_out;
  wire  regs_180_io_enable;
  wire  regs_181_clock;
  wire  regs_181_reset;
  wire [63:0] regs_181_io_in;
  wire [63:0] regs_181_io_init;
  wire [63:0] regs_181_io_out;
  wire  regs_181_io_enable;
  wire  regs_182_clock;
  wire  regs_182_reset;
  wire [63:0] regs_182_io_in;
  wire [63:0] regs_182_io_init;
  wire [63:0] regs_182_io_out;
  wire  regs_182_io_enable;
  wire  regs_183_clock;
  wire  regs_183_reset;
  wire [63:0] regs_183_io_in;
  wire [63:0] regs_183_io_init;
  wire [63:0] regs_183_io_out;
  wire  regs_183_io_enable;
  wire  regs_184_clock;
  wire  regs_184_reset;
  wire [63:0] regs_184_io_in;
  wire [63:0] regs_184_io_init;
  wire [63:0] regs_184_io_out;
  wire  regs_184_io_enable;
  wire  regs_185_clock;
  wire  regs_185_reset;
  wire [63:0] regs_185_io_in;
  wire [63:0] regs_185_io_init;
  wire [63:0] regs_185_io_out;
  wire  regs_185_io_enable;
  wire  regs_186_clock;
  wire  regs_186_reset;
  wire [63:0] regs_186_io_in;
  wire [63:0] regs_186_io_init;
  wire [63:0] regs_186_io_out;
  wire  regs_186_io_enable;
  wire  regs_187_clock;
  wire  regs_187_reset;
  wire [63:0] regs_187_io_in;
  wire [63:0] regs_187_io_init;
  wire [63:0] regs_187_io_out;
  wire  regs_187_io_enable;
  wire  regs_188_clock;
  wire  regs_188_reset;
  wire [63:0] regs_188_io_in;
  wire [63:0] regs_188_io_init;
  wire [63:0] regs_188_io_out;
  wire  regs_188_io_enable;
  wire  regs_189_clock;
  wire  regs_189_reset;
  wire [63:0] regs_189_io_in;
  wire [63:0] regs_189_io_init;
  wire [63:0] regs_189_io_out;
  wire  regs_189_io_enable;
  wire  regs_190_clock;
  wire  regs_190_reset;
  wire [63:0] regs_190_io_in;
  wire [63:0] regs_190_io_init;
  wire [63:0] regs_190_io_out;
  wire  regs_190_io_enable;
  wire  regs_191_clock;
  wire  regs_191_reset;
  wire [63:0] regs_191_io_in;
  wire [63:0] regs_191_io_init;
  wire [63:0] regs_191_io_out;
  wire  regs_191_io_enable;
  wire  regs_192_clock;
  wire  regs_192_reset;
  wire [63:0] regs_192_io_in;
  wire [63:0] regs_192_io_init;
  wire [63:0] regs_192_io_out;
  wire  regs_192_io_enable;
  wire  regs_193_clock;
  wire  regs_193_reset;
  wire [63:0] regs_193_io_in;
  wire [63:0] regs_193_io_init;
  wire [63:0] regs_193_io_out;
  wire  regs_193_io_enable;
  wire  regs_194_clock;
  wire  regs_194_reset;
  wire [63:0] regs_194_io_in;
  wire [63:0] regs_194_io_init;
  wire [63:0] regs_194_io_out;
  wire  regs_194_io_enable;
  wire  regs_195_clock;
  wire  regs_195_reset;
  wire [63:0] regs_195_io_in;
  wire [63:0] regs_195_io_init;
  wire [63:0] regs_195_io_out;
  wire  regs_195_io_enable;
  wire  regs_196_clock;
  wire  regs_196_reset;
  wire [63:0] regs_196_io_in;
  wire [63:0] regs_196_io_init;
  wire [63:0] regs_196_io_out;
  wire  regs_196_io_enable;
  wire  regs_197_clock;
  wire  regs_197_reset;
  wire [63:0] regs_197_io_in;
  wire [63:0] regs_197_io_init;
  wire [63:0] regs_197_io_out;
  wire  regs_197_io_enable;
  wire  regs_198_clock;
  wire  regs_198_reset;
  wire [63:0] regs_198_io_in;
  wire [63:0] regs_198_io_init;
  wire [63:0] regs_198_io_out;
  wire  regs_198_io_enable;
  wire  regs_199_clock;
  wire  regs_199_reset;
  wire [63:0] regs_199_io_in;
  wire [63:0] regs_199_io_init;
  wire [63:0] regs_199_io_out;
  wire  regs_199_io_enable;
  wire  regs_200_clock;
  wire  regs_200_reset;
  wire [63:0] regs_200_io_in;
  wire [63:0] regs_200_io_init;
  wire [63:0] regs_200_io_out;
  wire  regs_200_io_enable;
  wire  regs_201_clock;
  wire  regs_201_reset;
  wire [63:0] regs_201_io_in;
  wire [63:0] regs_201_io_init;
  wire [63:0] regs_201_io_out;
  wire  regs_201_io_enable;
  wire  regs_202_clock;
  wire  regs_202_reset;
  wire [63:0] regs_202_io_in;
  wire [63:0] regs_202_io_init;
  wire [63:0] regs_202_io_out;
  wire  regs_202_io_enable;
  wire  regs_203_clock;
  wire  regs_203_reset;
  wire [63:0] regs_203_io_in;
  wire [63:0] regs_203_io_init;
  wire [63:0] regs_203_io_out;
  wire  regs_203_io_enable;
  wire  regs_204_clock;
  wire  regs_204_reset;
  wire [63:0] regs_204_io_in;
  wire [63:0] regs_204_io_init;
  wire [63:0] regs_204_io_out;
  wire  regs_204_io_enable;
  wire  regs_205_clock;
  wire  regs_205_reset;
  wire [63:0] regs_205_io_in;
  wire [63:0] regs_205_io_init;
  wire [63:0] regs_205_io_out;
  wire  regs_205_io_enable;
  wire  regs_206_clock;
  wire  regs_206_reset;
  wire [63:0] regs_206_io_in;
  wire [63:0] regs_206_io_init;
  wire [63:0] regs_206_io_out;
  wire  regs_206_io_enable;
  wire  regs_207_clock;
  wire  regs_207_reset;
  wire [63:0] regs_207_io_in;
  wire [63:0] regs_207_io_init;
  wire [63:0] regs_207_io_out;
  wire  regs_207_io_enable;
  wire  regs_208_clock;
  wire  regs_208_reset;
  wire [63:0] regs_208_io_in;
  wire [63:0] regs_208_io_init;
  wire [63:0] regs_208_io_out;
  wire  regs_208_io_enable;
  wire  regs_209_clock;
  wire  regs_209_reset;
  wire [63:0] regs_209_io_in;
  wire [63:0] regs_209_io_init;
  wire [63:0] regs_209_io_out;
  wire  regs_209_io_enable;
  wire  regs_210_clock;
  wire  regs_210_reset;
  wire [63:0] regs_210_io_in;
  wire [63:0] regs_210_io_init;
  wire [63:0] regs_210_io_out;
  wire  regs_210_io_enable;
  wire  regs_211_clock;
  wire  regs_211_reset;
  wire [63:0] regs_211_io_in;
  wire [63:0] regs_211_io_init;
  wire [63:0] regs_211_io_out;
  wire  regs_211_io_enable;
  wire  regs_212_clock;
  wire  regs_212_reset;
  wire [63:0] regs_212_io_in;
  wire [63:0] regs_212_io_init;
  wire [63:0] regs_212_io_out;
  wire  regs_212_io_enable;
  wire  regs_213_clock;
  wire  regs_213_reset;
  wire [63:0] regs_213_io_in;
  wire [63:0] regs_213_io_init;
  wire [63:0] regs_213_io_out;
  wire  regs_213_io_enable;
  wire  regs_214_clock;
  wire  regs_214_reset;
  wire [63:0] regs_214_io_in;
  wire [63:0] regs_214_io_init;
  wire [63:0] regs_214_io_out;
  wire  regs_214_io_enable;
  wire  regs_215_clock;
  wire  regs_215_reset;
  wire [63:0] regs_215_io_in;
  wire [63:0] regs_215_io_init;
  wire [63:0] regs_215_io_out;
  wire  regs_215_io_enable;
  wire  regs_216_clock;
  wire  regs_216_reset;
  wire [63:0] regs_216_io_in;
  wire [63:0] regs_216_io_init;
  wire [63:0] regs_216_io_out;
  wire  regs_216_io_enable;
  wire  regs_217_clock;
  wire  regs_217_reset;
  wire [63:0] regs_217_io_in;
  wire [63:0] regs_217_io_init;
  wire [63:0] regs_217_io_out;
  wire  regs_217_io_enable;
  wire  regs_218_clock;
  wire  regs_218_reset;
  wire [63:0] regs_218_io_in;
  wire [63:0] regs_218_io_init;
  wire [63:0] regs_218_io_out;
  wire  regs_218_io_enable;
  wire  regs_219_clock;
  wire  regs_219_reset;
  wire [63:0] regs_219_io_in;
  wire [63:0] regs_219_io_init;
  wire [63:0] regs_219_io_out;
  wire  regs_219_io_enable;
  wire  regs_220_clock;
  wire  regs_220_reset;
  wire [63:0] regs_220_io_in;
  wire [63:0] regs_220_io_init;
  wire [63:0] regs_220_io_out;
  wire  regs_220_io_enable;
  wire  regs_221_clock;
  wire  regs_221_reset;
  wire [63:0] regs_221_io_in;
  wire [63:0] regs_221_io_init;
  wire [63:0] regs_221_io_out;
  wire  regs_221_io_enable;
  wire  regs_222_clock;
  wire  regs_222_reset;
  wire [63:0] regs_222_io_in;
  wire [63:0] regs_222_io_init;
  wire [63:0] regs_222_io_out;
  wire  regs_222_io_enable;
  wire  regs_223_clock;
  wire  regs_223_reset;
  wire [63:0] regs_223_io_in;
  wire [63:0] regs_223_io_init;
  wire [63:0] regs_223_io_out;
  wire  regs_223_io_enable;
  wire  regs_224_clock;
  wire  regs_224_reset;
  wire [63:0] regs_224_io_in;
  wire [63:0] regs_224_io_init;
  wire [63:0] regs_224_io_out;
  wire  regs_224_io_enable;
  wire  regs_225_clock;
  wire  regs_225_reset;
  wire [63:0] regs_225_io_in;
  wire [63:0] regs_225_io_init;
  wire [63:0] regs_225_io_out;
  wire  regs_225_io_enable;
  wire  regs_226_clock;
  wire  regs_226_reset;
  wire [63:0] regs_226_io_in;
  wire [63:0] regs_226_io_init;
  wire [63:0] regs_226_io_out;
  wire  regs_226_io_enable;
  wire  regs_227_clock;
  wire  regs_227_reset;
  wire [63:0] regs_227_io_in;
  wire [63:0] regs_227_io_init;
  wire [63:0] regs_227_io_out;
  wire  regs_227_io_enable;
  wire  regs_228_clock;
  wire  regs_228_reset;
  wire [63:0] regs_228_io_in;
  wire [63:0] regs_228_io_init;
  wire [63:0] regs_228_io_out;
  wire  regs_228_io_enable;
  wire  regs_229_clock;
  wire  regs_229_reset;
  wire [63:0] regs_229_io_in;
  wire [63:0] regs_229_io_init;
  wire [63:0] regs_229_io_out;
  wire  regs_229_io_enable;
  wire  regs_230_clock;
  wire  regs_230_reset;
  wire [63:0] regs_230_io_in;
  wire [63:0] regs_230_io_init;
  wire [63:0] regs_230_io_out;
  wire  regs_230_io_enable;
  wire  regs_231_clock;
  wire  regs_231_reset;
  wire [63:0] regs_231_io_in;
  wire [63:0] regs_231_io_init;
  wire [63:0] regs_231_io_out;
  wire  regs_231_io_enable;
  wire  regs_232_clock;
  wire  regs_232_reset;
  wire [63:0] regs_232_io_in;
  wire [63:0] regs_232_io_init;
  wire [63:0] regs_232_io_out;
  wire  regs_232_io_enable;
  wire  regs_233_clock;
  wire  regs_233_reset;
  wire [63:0] regs_233_io_in;
  wire [63:0] regs_233_io_init;
  wire [63:0] regs_233_io_out;
  wire  regs_233_io_enable;
  wire  regs_234_clock;
  wire  regs_234_reset;
  wire [63:0] regs_234_io_in;
  wire [63:0] regs_234_io_init;
  wire [63:0] regs_234_io_out;
  wire  regs_234_io_enable;
  wire  regs_235_clock;
  wire  regs_235_reset;
  wire [63:0] regs_235_io_in;
  wire [63:0] regs_235_io_init;
  wire [63:0] regs_235_io_out;
  wire  regs_235_io_enable;
  wire  regs_236_clock;
  wire  regs_236_reset;
  wire [63:0] regs_236_io_in;
  wire [63:0] regs_236_io_init;
  wire [63:0] regs_236_io_out;
  wire  regs_236_io_enable;
  wire  regs_237_clock;
  wire  regs_237_reset;
  wire [63:0] regs_237_io_in;
  wire [63:0] regs_237_io_init;
  wire [63:0] regs_237_io_out;
  wire  regs_237_io_enable;
  wire  regs_238_clock;
  wire  regs_238_reset;
  wire [63:0] regs_238_io_in;
  wire [63:0] regs_238_io_init;
  wire [63:0] regs_238_io_out;
  wire  regs_238_io_enable;
  wire  regs_239_clock;
  wire  regs_239_reset;
  wire [63:0] regs_239_io_in;
  wire [63:0] regs_239_io_init;
  wire [63:0] regs_239_io_out;
  wire  regs_239_io_enable;
  wire  regs_240_clock;
  wire  regs_240_reset;
  wire [63:0] regs_240_io_in;
  wire [63:0] regs_240_io_init;
  wire [63:0] regs_240_io_out;
  wire  regs_240_io_enable;
  wire  regs_241_clock;
  wire  regs_241_reset;
  wire [63:0] regs_241_io_in;
  wire [63:0] regs_241_io_init;
  wire [63:0] regs_241_io_out;
  wire  regs_241_io_enable;
  wire  regs_242_clock;
  wire  regs_242_reset;
  wire [63:0] regs_242_io_in;
  wire [63:0] regs_242_io_init;
  wire [63:0] regs_242_io_out;
  wire  regs_242_io_enable;
  wire  regs_243_clock;
  wire  regs_243_reset;
  wire [63:0] regs_243_io_in;
  wire [63:0] regs_243_io_init;
  wire [63:0] regs_243_io_out;
  wire  regs_243_io_enable;
  wire  regs_244_clock;
  wire  regs_244_reset;
  wire [63:0] regs_244_io_in;
  wire [63:0] regs_244_io_init;
  wire [63:0] regs_244_io_out;
  wire  regs_244_io_enable;
  wire  regs_245_clock;
  wire  regs_245_reset;
  wire [63:0] regs_245_io_in;
  wire [63:0] regs_245_io_init;
  wire [63:0] regs_245_io_out;
  wire  regs_245_io_enable;
  wire  regs_246_clock;
  wire  regs_246_reset;
  wire [63:0] regs_246_io_in;
  wire [63:0] regs_246_io_init;
  wire [63:0] regs_246_io_out;
  wire  regs_246_io_enable;
  wire  regs_247_clock;
  wire  regs_247_reset;
  wire [63:0] regs_247_io_in;
  wire [63:0] regs_247_io_init;
  wire [63:0] regs_247_io_out;
  wire  regs_247_io_enable;
  wire  regs_248_clock;
  wire  regs_248_reset;
  wire [63:0] regs_248_io_in;
  wire [63:0] regs_248_io_init;
  wire [63:0] regs_248_io_out;
  wire  regs_248_io_enable;
  wire  regs_249_clock;
  wire  regs_249_reset;
  wire [63:0] regs_249_io_in;
  wire [63:0] regs_249_io_init;
  wire [63:0] regs_249_io_out;
  wire  regs_249_io_enable;
  wire  regs_250_clock;
  wire  regs_250_reset;
  wire [63:0] regs_250_io_in;
  wire [63:0] regs_250_io_init;
  wire [63:0] regs_250_io_out;
  wire  regs_250_io_enable;
  wire  regs_251_clock;
  wire  regs_251_reset;
  wire [63:0] regs_251_io_in;
  wire [63:0] regs_251_io_init;
  wire [63:0] regs_251_io_out;
  wire  regs_251_io_enable;
  wire  regs_252_clock;
  wire  regs_252_reset;
  wire [63:0] regs_252_io_in;
  wire [63:0] regs_252_io_init;
  wire [63:0] regs_252_io_out;
  wire  regs_252_io_enable;
  wire  regs_253_clock;
  wire  regs_253_reset;
  wire [63:0] regs_253_io_in;
  wire [63:0] regs_253_io_init;
  wire [63:0] regs_253_io_out;
  wire  regs_253_io_enable;
  wire  regs_254_clock;
  wire  regs_254_reset;
  wire [63:0] regs_254_io_in;
  wire [63:0] regs_254_io_init;
  wire [63:0] regs_254_io_out;
  wire  regs_254_io_enable;
  wire  regs_255_clock;
  wire  regs_255_reset;
  wire [63:0] regs_255_io_in;
  wire [63:0] regs_255_io_init;
  wire [63:0] regs_255_io_out;
  wire  regs_255_io_enable;
  wire  regs_256_clock;
  wire  regs_256_reset;
  wire [63:0] regs_256_io_in;
  wire [63:0] regs_256_io_init;
  wire [63:0] regs_256_io_out;
  wire  regs_256_io_enable;
  wire  regs_257_clock;
  wire  regs_257_reset;
  wire [63:0] regs_257_io_in;
  wire [63:0] regs_257_io_init;
  wire [63:0] regs_257_io_out;
  wire  regs_257_io_enable;
  wire  regs_258_clock;
  wire  regs_258_reset;
  wire [63:0] regs_258_io_in;
  wire [63:0] regs_258_io_init;
  wire [63:0] regs_258_io_out;
  wire  regs_258_io_enable;
  wire  regs_259_clock;
  wire  regs_259_reset;
  wire [63:0] regs_259_io_in;
  wire [63:0] regs_259_io_init;
  wire [63:0] regs_259_io_out;
  wire  regs_259_io_enable;
  wire  regs_260_clock;
  wire  regs_260_reset;
  wire [63:0] regs_260_io_in;
  wire [63:0] regs_260_io_init;
  wire [63:0] regs_260_io_out;
  wire  regs_260_io_enable;
  wire  regs_261_clock;
  wire  regs_261_reset;
  wire [63:0] regs_261_io_in;
  wire [63:0] regs_261_io_init;
  wire [63:0] regs_261_io_out;
  wire  regs_261_io_enable;
  wire  regs_262_clock;
  wire  regs_262_reset;
  wire [63:0] regs_262_io_in;
  wire [63:0] regs_262_io_init;
  wire [63:0] regs_262_io_out;
  wire  regs_262_io_enable;
  wire  regs_263_clock;
  wire  regs_263_reset;
  wire [63:0] regs_263_io_in;
  wire [63:0] regs_263_io_init;
  wire [63:0] regs_263_io_out;
  wire  regs_263_io_enable;
  wire  regs_264_clock;
  wire  regs_264_reset;
  wire [63:0] regs_264_io_in;
  wire [63:0] regs_264_io_init;
  wire [63:0] regs_264_io_out;
  wire  regs_264_io_enable;
  wire  regs_265_clock;
  wire  regs_265_reset;
  wire [63:0] regs_265_io_in;
  wire [63:0] regs_265_io_init;
  wire [63:0] regs_265_io_out;
  wire  regs_265_io_enable;
  wire  regs_266_clock;
  wire  regs_266_reset;
  wire [63:0] regs_266_io_in;
  wire [63:0] regs_266_io_init;
  wire [63:0] regs_266_io_out;
  wire  regs_266_io_enable;
  wire  regs_267_clock;
  wire  regs_267_reset;
  wire [63:0] regs_267_io_in;
  wire [63:0] regs_267_io_init;
  wire [63:0] regs_267_io_out;
  wire  regs_267_io_enable;
  wire  regs_268_clock;
  wire  regs_268_reset;
  wire [63:0] regs_268_io_in;
  wire [63:0] regs_268_io_init;
  wire [63:0] regs_268_io_out;
  wire  regs_268_io_enable;
  wire  regs_269_clock;
  wire  regs_269_reset;
  wire [63:0] regs_269_io_in;
  wire [63:0] regs_269_io_init;
  wire [63:0] regs_269_io_out;
  wire  regs_269_io_enable;
  wire  regs_270_clock;
  wire  regs_270_reset;
  wire [63:0] regs_270_io_in;
  wire [63:0] regs_270_io_init;
  wire [63:0] regs_270_io_out;
  wire  regs_270_io_enable;
  wire  regs_271_clock;
  wire  regs_271_reset;
  wire [63:0] regs_271_io_in;
  wire [63:0] regs_271_io_init;
  wire [63:0] regs_271_io_out;
  wire  regs_271_io_enable;
  wire  regs_272_clock;
  wire  regs_272_reset;
  wire [63:0] regs_272_io_in;
  wire [63:0] regs_272_io_init;
  wire [63:0] regs_272_io_out;
  wire  regs_272_io_enable;
  wire  regs_273_clock;
  wire  regs_273_reset;
  wire [63:0] regs_273_io_in;
  wire [63:0] regs_273_io_init;
  wire [63:0] regs_273_io_out;
  wire  regs_273_io_enable;
  wire  regs_274_clock;
  wire  regs_274_reset;
  wire [63:0] regs_274_io_in;
  wire [63:0] regs_274_io_init;
  wire [63:0] regs_274_io_out;
  wire  regs_274_io_enable;
  wire  regs_275_clock;
  wire  regs_275_reset;
  wire [63:0] regs_275_io_in;
  wire [63:0] regs_275_io_init;
  wire [63:0] regs_275_io_out;
  wire  regs_275_io_enable;
  wire  regs_276_clock;
  wire  regs_276_reset;
  wire [63:0] regs_276_io_in;
  wire [63:0] regs_276_io_init;
  wire [63:0] regs_276_io_out;
  wire  regs_276_io_enable;
  wire  regs_277_clock;
  wire  regs_277_reset;
  wire [63:0] regs_277_io_in;
  wire [63:0] regs_277_io_init;
  wire [63:0] regs_277_io_out;
  wire  regs_277_io_enable;
  wire  regs_278_clock;
  wire  regs_278_reset;
  wire [63:0] regs_278_io_in;
  wire [63:0] regs_278_io_init;
  wire [63:0] regs_278_io_out;
  wire  regs_278_io_enable;
  wire  regs_279_clock;
  wire  regs_279_reset;
  wire [63:0] regs_279_io_in;
  wire [63:0] regs_279_io_init;
  wire [63:0] regs_279_io_out;
  wire  regs_279_io_enable;
  wire  regs_280_clock;
  wire  regs_280_reset;
  wire [63:0] regs_280_io_in;
  wire [63:0] regs_280_io_init;
  wire [63:0] regs_280_io_out;
  wire  regs_280_io_enable;
  wire  regs_281_clock;
  wire  regs_281_reset;
  wire [63:0] regs_281_io_in;
  wire [63:0] regs_281_io_init;
  wire [63:0] regs_281_io_out;
  wire  regs_281_io_enable;
  wire  regs_282_clock;
  wire  regs_282_reset;
  wire [63:0] regs_282_io_in;
  wire [63:0] regs_282_io_init;
  wire [63:0] regs_282_io_out;
  wire  regs_282_io_enable;
  wire  regs_283_clock;
  wire  regs_283_reset;
  wire [63:0] regs_283_io_in;
  wire [63:0] regs_283_io_init;
  wire [63:0] regs_283_io_out;
  wire  regs_283_io_enable;
  wire  regs_284_clock;
  wire  regs_284_reset;
  wire [63:0] regs_284_io_in;
  wire [63:0] regs_284_io_init;
  wire [63:0] regs_284_io_out;
  wire  regs_284_io_enable;
  wire  regs_285_clock;
  wire  regs_285_reset;
  wire [63:0] regs_285_io_in;
  wire [63:0] regs_285_io_init;
  wire [63:0] regs_285_io_out;
  wire  regs_285_io_enable;
  wire  regs_286_clock;
  wire  regs_286_reset;
  wire [63:0] regs_286_io_in;
  wire [63:0] regs_286_io_init;
  wire [63:0] regs_286_io_out;
  wire  regs_286_io_enable;
  wire  regs_287_clock;
  wire  regs_287_reset;
  wire [63:0] regs_287_io_in;
  wire [63:0] regs_287_io_init;
  wire [63:0] regs_287_io_out;
  wire  regs_287_io_enable;
  wire  regs_288_clock;
  wire  regs_288_reset;
  wire [63:0] regs_288_io_in;
  wire [63:0] regs_288_io_init;
  wire [63:0] regs_288_io_out;
  wire  regs_288_io_enable;
  wire  regs_289_clock;
  wire  regs_289_reset;
  wire [63:0] regs_289_io_in;
  wire [63:0] regs_289_io_init;
  wire [63:0] regs_289_io_out;
  wire  regs_289_io_enable;
  wire  regs_290_clock;
  wire  regs_290_reset;
  wire [63:0] regs_290_io_in;
  wire [63:0] regs_290_io_init;
  wire [63:0] regs_290_io_out;
  wire  regs_290_io_enable;
  wire  regs_291_clock;
  wire  regs_291_reset;
  wire [63:0] regs_291_io_in;
  wire [63:0] regs_291_io_init;
  wire [63:0] regs_291_io_out;
  wire  regs_291_io_enable;
  wire  regs_292_clock;
  wire  regs_292_reset;
  wire [63:0] regs_292_io_in;
  wire [63:0] regs_292_io_init;
  wire [63:0] regs_292_io_out;
  wire  regs_292_io_enable;
  wire  regs_293_clock;
  wire  regs_293_reset;
  wire [63:0] regs_293_io_in;
  wire [63:0] regs_293_io_init;
  wire [63:0] regs_293_io_out;
  wire  regs_293_io_enable;
  wire  regs_294_clock;
  wire  regs_294_reset;
  wire [63:0] regs_294_io_in;
  wire [63:0] regs_294_io_init;
  wire [63:0] regs_294_io_out;
  wire  regs_294_io_enable;
  wire  regs_295_clock;
  wire  regs_295_reset;
  wire [63:0] regs_295_io_in;
  wire [63:0] regs_295_io_init;
  wire [63:0] regs_295_io_out;
  wire  regs_295_io_enable;
  wire  regs_296_clock;
  wire  regs_296_reset;
  wire [63:0] regs_296_io_in;
  wire [63:0] regs_296_io_init;
  wire [63:0] regs_296_io_out;
  wire  regs_296_io_enable;
  wire  regs_297_clock;
  wire  regs_297_reset;
  wire [63:0] regs_297_io_in;
  wire [63:0] regs_297_io_init;
  wire [63:0] regs_297_io_out;
  wire  regs_297_io_enable;
  wire  regs_298_clock;
  wire  regs_298_reset;
  wire [63:0] regs_298_io_in;
  wire [63:0] regs_298_io_init;
  wire [63:0] regs_298_io_out;
  wire  regs_298_io_enable;
  wire  regs_299_clock;
  wire  regs_299_reset;
  wire [63:0] regs_299_io_in;
  wire [63:0] regs_299_io_init;
  wire [63:0] regs_299_io_out;
  wire  regs_299_io_enable;
  wire  regs_300_clock;
  wire  regs_300_reset;
  wire [63:0] regs_300_io_in;
  wire [63:0] regs_300_io_init;
  wire [63:0] regs_300_io_out;
  wire  regs_300_io_enable;
  wire  regs_301_clock;
  wire  regs_301_reset;
  wire [63:0] regs_301_io_in;
  wire [63:0] regs_301_io_init;
  wire [63:0] regs_301_io_out;
  wire  regs_301_io_enable;
  wire  regs_302_clock;
  wire  regs_302_reset;
  wire [63:0] regs_302_io_in;
  wire [63:0] regs_302_io_init;
  wire [63:0] regs_302_io_out;
  wire  regs_302_io_enable;
  wire  regs_303_clock;
  wire  regs_303_reset;
  wire [63:0] regs_303_io_in;
  wire [63:0] regs_303_io_init;
  wire [63:0] regs_303_io_out;
  wire  regs_303_io_enable;
  wire  regs_304_clock;
  wire  regs_304_reset;
  wire [63:0] regs_304_io_in;
  wire [63:0] regs_304_io_init;
  wire [63:0] regs_304_io_out;
  wire  regs_304_io_enable;
  wire  regs_305_clock;
  wire  regs_305_reset;
  wire [63:0] regs_305_io_in;
  wire [63:0] regs_305_io_init;
  wire [63:0] regs_305_io_out;
  wire  regs_305_io_enable;
  wire  regs_306_clock;
  wire  regs_306_reset;
  wire [63:0] regs_306_io_in;
  wire [63:0] regs_306_io_init;
  wire [63:0] regs_306_io_out;
  wire  regs_306_io_enable;
  wire  regs_307_clock;
  wire  regs_307_reset;
  wire [63:0] regs_307_io_in;
  wire [63:0] regs_307_io_init;
  wire [63:0] regs_307_io_out;
  wire  regs_307_io_enable;
  wire  regs_308_clock;
  wire  regs_308_reset;
  wire [63:0] regs_308_io_in;
  wire [63:0] regs_308_io_init;
  wire [63:0] regs_308_io_out;
  wire  regs_308_io_enable;
  wire  regs_309_clock;
  wire  regs_309_reset;
  wire [63:0] regs_309_io_in;
  wire [63:0] regs_309_io_init;
  wire [63:0] regs_309_io_out;
  wire  regs_309_io_enable;
  wire  regs_310_clock;
  wire  regs_310_reset;
  wire [63:0] regs_310_io_in;
  wire [63:0] regs_310_io_init;
  wire [63:0] regs_310_io_out;
  wire  regs_310_io_enable;
  wire  regs_311_clock;
  wire  regs_311_reset;
  wire [63:0] regs_311_io_in;
  wire [63:0] regs_311_io_init;
  wire [63:0] regs_311_io_out;
  wire  regs_311_io_enable;
  wire  regs_312_clock;
  wire  regs_312_reset;
  wire [63:0] regs_312_io_in;
  wire [63:0] regs_312_io_init;
  wire [63:0] regs_312_io_out;
  wire  regs_312_io_enable;
  wire  regs_313_clock;
  wire  regs_313_reset;
  wire [63:0] regs_313_io_in;
  wire [63:0] regs_313_io_init;
  wire [63:0] regs_313_io_out;
  wire  regs_313_io_enable;
  wire  regs_314_clock;
  wire  regs_314_reset;
  wire [63:0] regs_314_io_in;
  wire [63:0] regs_314_io_init;
  wire [63:0] regs_314_io_out;
  wire  regs_314_io_enable;
  wire  regs_315_clock;
  wire  regs_315_reset;
  wire [63:0] regs_315_io_in;
  wire [63:0] regs_315_io_init;
  wire [63:0] regs_315_io_out;
  wire  regs_315_io_enable;
  wire  regs_316_clock;
  wire  regs_316_reset;
  wire [63:0] regs_316_io_in;
  wire [63:0] regs_316_io_init;
  wire [63:0] regs_316_io_out;
  wire  regs_316_io_enable;
  wire  regs_317_clock;
  wire  regs_317_reset;
  wire [63:0] regs_317_io_in;
  wire [63:0] regs_317_io_init;
  wire [63:0] regs_317_io_out;
  wire  regs_317_io_enable;
  wire  regs_318_clock;
  wire  regs_318_reset;
  wire [63:0] regs_318_io_in;
  wire [63:0] regs_318_io_init;
  wire [63:0] regs_318_io_out;
  wire  regs_318_io_enable;
  wire  regs_319_clock;
  wire  regs_319_reset;
  wire [63:0] regs_319_io_in;
  wire [63:0] regs_319_io_init;
  wire [63:0] regs_319_io_out;
  wire  regs_319_io_enable;
  wire  regs_320_clock;
  wire  regs_320_reset;
  wire [63:0] regs_320_io_in;
  wire [63:0] regs_320_io_init;
  wire [63:0] regs_320_io_out;
  wire  regs_320_io_enable;
  wire  regs_321_clock;
  wire  regs_321_reset;
  wire [63:0] regs_321_io_in;
  wire [63:0] regs_321_io_init;
  wire [63:0] regs_321_io_out;
  wire  regs_321_io_enable;
  wire  regs_322_clock;
  wire  regs_322_reset;
  wire [63:0] regs_322_io_in;
  wire [63:0] regs_322_io_init;
  wire [63:0] regs_322_io_out;
  wire  regs_322_io_enable;
  wire  regs_323_clock;
  wire  regs_323_reset;
  wire [63:0] regs_323_io_in;
  wire [63:0] regs_323_io_init;
  wire [63:0] regs_323_io_out;
  wire  regs_323_io_enable;
  wire  regs_324_clock;
  wire  regs_324_reset;
  wire [63:0] regs_324_io_in;
  wire [63:0] regs_324_io_init;
  wire [63:0] regs_324_io_out;
  wire  regs_324_io_enable;
  wire  regs_325_clock;
  wire  regs_325_reset;
  wire [63:0] regs_325_io_in;
  wire [63:0] regs_325_io_init;
  wire [63:0] regs_325_io_out;
  wire  regs_325_io_enable;
  wire  regs_326_clock;
  wire  regs_326_reset;
  wire [63:0] regs_326_io_in;
  wire [63:0] regs_326_io_init;
  wire [63:0] regs_326_io_out;
  wire  regs_326_io_enable;
  wire  regs_327_clock;
  wire  regs_327_reset;
  wire [63:0] regs_327_io_in;
  wire [63:0] regs_327_io_init;
  wire [63:0] regs_327_io_out;
  wire  regs_327_io_enable;
  wire  regs_328_clock;
  wire  regs_328_reset;
  wire [63:0] regs_328_io_in;
  wire [63:0] regs_328_io_init;
  wire [63:0] regs_328_io_out;
  wire  regs_328_io_enable;
  wire  regs_329_clock;
  wire  regs_329_reset;
  wire [63:0] regs_329_io_in;
  wire [63:0] regs_329_io_init;
  wire [63:0] regs_329_io_out;
  wire  regs_329_io_enable;
  wire  regs_330_clock;
  wire  regs_330_reset;
  wire [63:0] regs_330_io_in;
  wire [63:0] regs_330_io_init;
  wire [63:0] regs_330_io_out;
  wire  regs_330_io_enable;
  wire  regs_331_clock;
  wire  regs_331_reset;
  wire [63:0] regs_331_io_in;
  wire [63:0] regs_331_io_init;
  wire [63:0] regs_331_io_out;
  wire  regs_331_io_enable;
  wire  regs_332_clock;
  wire  regs_332_reset;
  wire [63:0] regs_332_io_in;
  wire [63:0] regs_332_io_init;
  wire [63:0] regs_332_io_out;
  wire  regs_332_io_enable;
  wire  regs_333_clock;
  wire  regs_333_reset;
  wire [63:0] regs_333_io_in;
  wire [63:0] regs_333_io_init;
  wire [63:0] regs_333_io_out;
  wire  regs_333_io_enable;
  wire  regs_334_clock;
  wire  regs_334_reset;
  wire [63:0] regs_334_io_in;
  wire [63:0] regs_334_io_init;
  wire [63:0] regs_334_io_out;
  wire  regs_334_io_enable;
  wire  regs_335_clock;
  wire  regs_335_reset;
  wire [63:0] regs_335_io_in;
  wire [63:0] regs_335_io_init;
  wire [63:0] regs_335_io_out;
  wire  regs_335_io_enable;
  wire  regs_336_clock;
  wire  regs_336_reset;
  wire [63:0] regs_336_io_in;
  wire [63:0] regs_336_io_init;
  wire [63:0] regs_336_io_out;
  wire  regs_336_io_enable;
  wire  regs_337_clock;
  wire  regs_337_reset;
  wire [63:0] regs_337_io_in;
  wire [63:0] regs_337_io_init;
  wire [63:0] regs_337_io_out;
  wire  regs_337_io_enable;
  wire  regs_338_clock;
  wire  regs_338_reset;
  wire [63:0] regs_338_io_in;
  wire [63:0] regs_338_io_init;
  wire [63:0] regs_338_io_out;
  wire  regs_338_io_enable;
  wire  regs_339_clock;
  wire  regs_339_reset;
  wire [63:0] regs_339_io_in;
  wire [63:0] regs_339_io_init;
  wire [63:0] regs_339_io_out;
  wire  regs_339_io_enable;
  wire  regs_340_clock;
  wire  regs_340_reset;
  wire [63:0] regs_340_io_in;
  wire [63:0] regs_340_io_init;
  wire [63:0] regs_340_io_out;
  wire  regs_340_io_enable;
  wire  regs_341_clock;
  wire  regs_341_reset;
  wire [63:0] regs_341_io_in;
  wire [63:0] regs_341_io_init;
  wire [63:0] regs_341_io_out;
  wire  regs_341_io_enable;
  wire  regs_342_clock;
  wire  regs_342_reset;
  wire [63:0] regs_342_io_in;
  wire [63:0] regs_342_io_init;
  wire [63:0] regs_342_io_out;
  wire  regs_342_io_enable;
  wire  regs_343_clock;
  wire  regs_343_reset;
  wire [63:0] regs_343_io_in;
  wire [63:0] regs_343_io_init;
  wire [63:0] regs_343_io_out;
  wire  regs_343_io_enable;
  wire  regs_344_clock;
  wire  regs_344_reset;
  wire [63:0] regs_344_io_in;
  wire [63:0] regs_344_io_init;
  wire [63:0] regs_344_io_out;
  wire  regs_344_io_enable;
  wire  regs_345_clock;
  wire  regs_345_reset;
  wire [63:0] regs_345_io_in;
  wire [63:0] regs_345_io_init;
  wire [63:0] regs_345_io_out;
  wire  regs_345_io_enable;
  wire  regs_346_clock;
  wire  regs_346_reset;
  wire [63:0] regs_346_io_in;
  wire [63:0] regs_346_io_init;
  wire [63:0] regs_346_io_out;
  wire  regs_346_io_enable;
  wire  regs_347_clock;
  wire  regs_347_reset;
  wire [63:0] regs_347_io_in;
  wire [63:0] regs_347_io_init;
  wire [63:0] regs_347_io_out;
  wire  regs_347_io_enable;
  wire  regs_348_clock;
  wire  regs_348_reset;
  wire [63:0] regs_348_io_in;
  wire [63:0] regs_348_io_init;
  wire [63:0] regs_348_io_out;
  wire  regs_348_io_enable;
  wire  regs_349_clock;
  wire  regs_349_reset;
  wire [63:0] regs_349_io_in;
  wire [63:0] regs_349_io_init;
  wire [63:0] regs_349_io_out;
  wire  regs_349_io_enable;
  wire  regs_350_clock;
  wire  regs_350_reset;
  wire [63:0] regs_350_io_in;
  wire [63:0] regs_350_io_init;
  wire [63:0] regs_350_io_out;
  wire  regs_350_io_enable;
  wire  regs_351_clock;
  wire  regs_351_reset;
  wire [63:0] regs_351_io_in;
  wire [63:0] regs_351_io_init;
  wire [63:0] regs_351_io_out;
  wire  regs_351_io_enable;
  wire  regs_352_clock;
  wire  regs_352_reset;
  wire [63:0] regs_352_io_in;
  wire [63:0] regs_352_io_init;
  wire [63:0] regs_352_io_out;
  wire  regs_352_io_enable;
  wire  regs_353_clock;
  wire  regs_353_reset;
  wire [63:0] regs_353_io_in;
  wire [63:0] regs_353_io_init;
  wire [63:0] regs_353_io_out;
  wire  regs_353_io_enable;
  wire  regs_354_clock;
  wire  regs_354_reset;
  wire [63:0] regs_354_io_in;
  wire [63:0] regs_354_io_init;
  wire [63:0] regs_354_io_out;
  wire  regs_354_io_enable;
  wire  regs_355_clock;
  wire  regs_355_reset;
  wire [63:0] regs_355_io_in;
  wire [63:0] regs_355_io_init;
  wire [63:0] regs_355_io_out;
  wire  regs_355_io_enable;
  wire  regs_356_clock;
  wire  regs_356_reset;
  wire [63:0] regs_356_io_in;
  wire [63:0] regs_356_io_init;
  wire [63:0] regs_356_io_out;
  wire  regs_356_io_enable;
  wire  regs_357_clock;
  wire  regs_357_reset;
  wire [63:0] regs_357_io_in;
  wire [63:0] regs_357_io_init;
  wire [63:0] regs_357_io_out;
  wire  regs_357_io_enable;
  wire  regs_358_clock;
  wire  regs_358_reset;
  wire [63:0] regs_358_io_in;
  wire [63:0] regs_358_io_init;
  wire [63:0] regs_358_io_out;
  wire  regs_358_io_enable;
  wire  regs_359_clock;
  wire  regs_359_reset;
  wire [63:0] regs_359_io_in;
  wire [63:0] regs_359_io_init;
  wire [63:0] regs_359_io_out;
  wire  regs_359_io_enable;
  wire  regs_360_clock;
  wire  regs_360_reset;
  wire [63:0] regs_360_io_in;
  wire [63:0] regs_360_io_init;
  wire [63:0] regs_360_io_out;
  wire  regs_360_io_enable;
  wire  regs_361_clock;
  wire  regs_361_reset;
  wire [63:0] regs_361_io_in;
  wire [63:0] regs_361_io_init;
  wire [63:0] regs_361_io_out;
  wire  regs_361_io_enable;
  wire  regs_362_clock;
  wire  regs_362_reset;
  wire [63:0] regs_362_io_in;
  wire [63:0] regs_362_io_init;
  wire [63:0] regs_362_io_out;
  wire  regs_362_io_enable;
  wire  regs_363_clock;
  wire  regs_363_reset;
  wire [63:0] regs_363_io_in;
  wire [63:0] regs_363_io_init;
  wire [63:0] regs_363_io_out;
  wire  regs_363_io_enable;
  wire  regs_364_clock;
  wire  regs_364_reset;
  wire [63:0] regs_364_io_in;
  wire [63:0] regs_364_io_init;
  wire [63:0] regs_364_io_out;
  wire  regs_364_io_enable;
  wire  regs_365_clock;
  wire  regs_365_reset;
  wire [63:0] regs_365_io_in;
  wire [63:0] regs_365_io_init;
  wire [63:0] regs_365_io_out;
  wire  regs_365_io_enable;
  wire  regs_366_clock;
  wire  regs_366_reset;
  wire [63:0] regs_366_io_in;
  wire [63:0] regs_366_io_init;
  wire [63:0] regs_366_io_out;
  wire  regs_366_io_enable;
  wire  regs_367_clock;
  wire  regs_367_reset;
  wire [63:0] regs_367_io_in;
  wire [63:0] regs_367_io_init;
  wire [63:0] regs_367_io_out;
  wire  regs_367_io_enable;
  wire  regs_368_clock;
  wire  regs_368_reset;
  wire [63:0] regs_368_io_in;
  wire [63:0] regs_368_io_init;
  wire [63:0] regs_368_io_out;
  wire  regs_368_io_enable;
  wire  regs_369_clock;
  wire  regs_369_reset;
  wire [63:0] regs_369_io_in;
  wire [63:0] regs_369_io_init;
  wire [63:0] regs_369_io_out;
  wire  regs_369_io_enable;
  wire  regs_370_clock;
  wire  regs_370_reset;
  wire [63:0] regs_370_io_in;
  wire [63:0] regs_370_io_init;
  wire [63:0] regs_370_io_out;
  wire  regs_370_io_enable;
  wire  regs_371_clock;
  wire  regs_371_reset;
  wire [63:0] regs_371_io_in;
  wire [63:0] regs_371_io_init;
  wire [63:0] regs_371_io_out;
  wire  regs_371_io_enable;
  wire  regs_372_clock;
  wire  regs_372_reset;
  wire [63:0] regs_372_io_in;
  wire [63:0] regs_372_io_init;
  wire [63:0] regs_372_io_out;
  wire  regs_372_io_enable;
  wire  regs_373_clock;
  wire  regs_373_reset;
  wire [63:0] regs_373_io_in;
  wire [63:0] regs_373_io_init;
  wire [63:0] regs_373_io_out;
  wire  regs_373_io_enable;
  wire  regs_374_clock;
  wire  regs_374_reset;
  wire [63:0] regs_374_io_in;
  wire [63:0] regs_374_io_init;
  wire [63:0] regs_374_io_out;
  wire  regs_374_io_enable;
  wire  regs_375_clock;
  wire  regs_375_reset;
  wire [63:0] regs_375_io_in;
  wire [63:0] regs_375_io_init;
  wire [63:0] regs_375_io_out;
  wire  regs_375_io_enable;
  wire  regs_376_clock;
  wire  regs_376_reset;
  wire [63:0] regs_376_io_in;
  wire [63:0] regs_376_io_init;
  wire [63:0] regs_376_io_out;
  wire  regs_376_io_enable;
  wire  regs_377_clock;
  wire  regs_377_reset;
  wire [63:0] regs_377_io_in;
  wire [63:0] regs_377_io_init;
  wire [63:0] regs_377_io_out;
  wire  regs_377_io_enable;
  wire  regs_378_clock;
  wire  regs_378_reset;
  wire [63:0] regs_378_io_in;
  wire [63:0] regs_378_io_init;
  wire [63:0] regs_378_io_out;
  wire  regs_378_io_enable;
  wire  regs_379_clock;
  wire  regs_379_reset;
  wire [63:0] regs_379_io_in;
  wire [63:0] regs_379_io_init;
  wire [63:0] regs_379_io_out;
  wire  regs_379_io_enable;
  wire  regs_380_clock;
  wire  regs_380_reset;
  wire [63:0] regs_380_io_in;
  wire [63:0] regs_380_io_init;
  wire [63:0] regs_380_io_out;
  wire  regs_380_io_enable;
  wire  regs_381_clock;
  wire  regs_381_reset;
  wire [63:0] regs_381_io_in;
  wire [63:0] regs_381_io_init;
  wire [63:0] regs_381_io_out;
  wire  regs_381_io_enable;
  wire  regs_382_clock;
  wire  regs_382_reset;
  wire [63:0] regs_382_io_in;
  wire [63:0] regs_382_io_init;
  wire [63:0] regs_382_io_out;
  wire  regs_382_io_enable;
  wire  regs_383_clock;
  wire  regs_383_reset;
  wire [63:0] regs_383_io_in;
  wire [63:0] regs_383_io_init;
  wire [63:0] regs_383_io_out;
  wire  regs_383_io_enable;
  wire  regs_384_clock;
  wire  regs_384_reset;
  wire [63:0] regs_384_io_in;
  wire [63:0] regs_384_io_init;
  wire [63:0] regs_384_io_out;
  wire  regs_384_io_enable;
  wire  regs_385_clock;
  wire  regs_385_reset;
  wire [63:0] regs_385_io_in;
  wire [63:0] regs_385_io_init;
  wire [63:0] regs_385_io_out;
  wire  regs_385_io_enable;
  wire  regs_386_clock;
  wire  regs_386_reset;
  wire [63:0] regs_386_io_in;
  wire [63:0] regs_386_io_init;
  wire [63:0] regs_386_io_out;
  wire  regs_386_io_enable;
  wire  regs_387_clock;
  wire  regs_387_reset;
  wire [63:0] regs_387_io_in;
  wire [63:0] regs_387_io_init;
  wire [63:0] regs_387_io_out;
  wire  regs_387_io_enable;
  wire  regs_388_clock;
  wire  regs_388_reset;
  wire [63:0] regs_388_io_in;
  wire [63:0] regs_388_io_init;
  wire [63:0] regs_388_io_out;
  wire  regs_388_io_enable;
  wire  regs_389_clock;
  wire  regs_389_reset;
  wire [63:0] regs_389_io_in;
  wire [63:0] regs_389_io_init;
  wire [63:0] regs_389_io_out;
  wire  regs_389_io_enable;
  wire  regs_390_clock;
  wire  regs_390_reset;
  wire [63:0] regs_390_io_in;
  wire [63:0] regs_390_io_init;
  wire [63:0] regs_390_io_out;
  wire  regs_390_io_enable;
  wire  regs_391_clock;
  wire  regs_391_reset;
  wire [63:0] regs_391_io_in;
  wire [63:0] regs_391_io_init;
  wire [63:0] regs_391_io_out;
  wire  regs_391_io_enable;
  wire  regs_392_clock;
  wire  regs_392_reset;
  wire [63:0] regs_392_io_in;
  wire [63:0] regs_392_io_init;
  wire [63:0] regs_392_io_out;
  wire  regs_392_io_enable;
  wire  regs_393_clock;
  wire  regs_393_reset;
  wire [63:0] regs_393_io_in;
  wire [63:0] regs_393_io_init;
  wire [63:0] regs_393_io_out;
  wire  regs_393_io_enable;
  wire  regs_394_clock;
  wire  regs_394_reset;
  wire [63:0] regs_394_io_in;
  wire [63:0] regs_394_io_init;
  wire [63:0] regs_394_io_out;
  wire  regs_394_io_enable;
  wire  regs_395_clock;
  wire  regs_395_reset;
  wire [63:0] regs_395_io_in;
  wire [63:0] regs_395_io_init;
  wire [63:0] regs_395_io_out;
  wire  regs_395_io_enable;
  wire  regs_396_clock;
  wire  regs_396_reset;
  wire [63:0] regs_396_io_in;
  wire [63:0] regs_396_io_init;
  wire [63:0] regs_396_io_out;
  wire  regs_396_io_enable;
  wire  regs_397_clock;
  wire  regs_397_reset;
  wire [63:0] regs_397_io_in;
  wire [63:0] regs_397_io_init;
  wire [63:0] regs_397_io_out;
  wire  regs_397_io_enable;
  wire  regs_398_clock;
  wire  regs_398_reset;
  wire [63:0] regs_398_io_in;
  wire [63:0] regs_398_io_init;
  wire [63:0] regs_398_io_out;
  wire  regs_398_io_enable;
  wire  regs_399_clock;
  wire  regs_399_reset;
  wire [63:0] regs_399_io_in;
  wire [63:0] regs_399_io_init;
  wire [63:0] regs_399_io_out;
  wire  regs_399_io_enable;
  wire  regs_400_clock;
  wire  regs_400_reset;
  wire [63:0] regs_400_io_in;
  wire [63:0] regs_400_io_init;
  wire [63:0] regs_400_io_out;
  wire  regs_400_io_enable;
  wire  regs_401_clock;
  wire  regs_401_reset;
  wire [63:0] regs_401_io_in;
  wire [63:0] regs_401_io_init;
  wire [63:0] regs_401_io_out;
  wire  regs_401_io_enable;
  wire  regs_402_clock;
  wire  regs_402_reset;
  wire [63:0] regs_402_io_in;
  wire [63:0] regs_402_io_init;
  wire [63:0] regs_402_io_out;
  wire  regs_402_io_enable;
  wire  regs_403_clock;
  wire  regs_403_reset;
  wire [63:0] regs_403_io_in;
  wire [63:0] regs_403_io_init;
  wire [63:0] regs_403_io_out;
  wire  regs_403_io_enable;
  wire  regs_404_clock;
  wire  regs_404_reset;
  wire [63:0] regs_404_io_in;
  wire [63:0] regs_404_io_init;
  wire [63:0] regs_404_io_out;
  wire  regs_404_io_enable;
  wire  regs_405_clock;
  wire  regs_405_reset;
  wire [63:0] regs_405_io_in;
  wire [63:0] regs_405_io_init;
  wire [63:0] regs_405_io_out;
  wire  regs_405_io_enable;
  wire  regs_406_clock;
  wire  regs_406_reset;
  wire [63:0] regs_406_io_in;
  wire [63:0] regs_406_io_init;
  wire [63:0] regs_406_io_out;
  wire  regs_406_io_enable;
  wire  regs_407_clock;
  wire  regs_407_reset;
  wire [63:0] regs_407_io_in;
  wire [63:0] regs_407_io_init;
  wire [63:0] regs_407_io_out;
  wire  regs_407_io_enable;
  wire  regs_408_clock;
  wire  regs_408_reset;
  wire [63:0] regs_408_io_in;
  wire [63:0] regs_408_io_init;
  wire [63:0] regs_408_io_out;
  wire  regs_408_io_enable;
  wire  regs_409_clock;
  wire  regs_409_reset;
  wire [63:0] regs_409_io_in;
  wire [63:0] regs_409_io_init;
  wire [63:0] regs_409_io_out;
  wire  regs_409_io_enable;
  wire  regs_410_clock;
  wire  regs_410_reset;
  wire [63:0] regs_410_io_in;
  wire [63:0] regs_410_io_init;
  wire [63:0] regs_410_io_out;
  wire  regs_410_io_enable;
  wire  regs_411_clock;
  wire  regs_411_reset;
  wire [63:0] regs_411_io_in;
  wire [63:0] regs_411_io_init;
  wire [63:0] regs_411_io_out;
  wire  regs_411_io_enable;
  wire  regs_412_clock;
  wire  regs_412_reset;
  wire [63:0] regs_412_io_in;
  wire [63:0] regs_412_io_init;
  wire [63:0] regs_412_io_out;
  wire  regs_412_io_enable;
  wire  regs_413_clock;
  wire  regs_413_reset;
  wire [63:0] regs_413_io_in;
  wire [63:0] regs_413_io_init;
  wire [63:0] regs_413_io_out;
  wire  regs_413_io_enable;
  wire  regs_414_clock;
  wire  regs_414_reset;
  wire [63:0] regs_414_io_in;
  wire [63:0] regs_414_io_init;
  wire [63:0] regs_414_io_out;
  wire  regs_414_io_enable;
  wire  regs_415_clock;
  wire  regs_415_reset;
  wire [63:0] regs_415_io_in;
  wire [63:0] regs_415_io_init;
  wire [63:0] regs_415_io_out;
  wire  regs_415_io_enable;
  wire  regs_416_clock;
  wire  regs_416_reset;
  wire [63:0] regs_416_io_in;
  wire [63:0] regs_416_io_init;
  wire [63:0] regs_416_io_out;
  wire  regs_416_io_enable;
  wire  regs_417_clock;
  wire  regs_417_reset;
  wire [63:0] regs_417_io_in;
  wire [63:0] regs_417_io_init;
  wire [63:0] regs_417_io_out;
  wire  regs_417_io_enable;
  wire  regs_418_clock;
  wire  regs_418_reset;
  wire [63:0] regs_418_io_in;
  wire [63:0] regs_418_io_init;
  wire [63:0] regs_418_io_out;
  wire  regs_418_io_enable;
  wire  regs_419_clock;
  wire  regs_419_reset;
  wire [63:0] regs_419_io_in;
  wire [63:0] regs_419_io_init;
  wire [63:0] regs_419_io_out;
  wire  regs_419_io_enable;
  wire  regs_420_clock;
  wire  regs_420_reset;
  wire [63:0] regs_420_io_in;
  wire [63:0] regs_420_io_init;
  wire [63:0] regs_420_io_out;
  wire  regs_420_io_enable;
  wire  regs_421_clock;
  wire  regs_421_reset;
  wire [63:0] regs_421_io_in;
  wire [63:0] regs_421_io_init;
  wire [63:0] regs_421_io_out;
  wire  regs_421_io_enable;
  wire  regs_422_clock;
  wire  regs_422_reset;
  wire [63:0] regs_422_io_in;
  wire [63:0] regs_422_io_init;
  wire [63:0] regs_422_io_out;
  wire  regs_422_io_enable;
  wire  regs_423_clock;
  wire  regs_423_reset;
  wire [63:0] regs_423_io_in;
  wire [63:0] regs_423_io_init;
  wire [63:0] regs_423_io_out;
  wire  regs_423_io_enable;
  wire  regs_424_clock;
  wire  regs_424_reset;
  wire [63:0] regs_424_io_in;
  wire [63:0] regs_424_io_init;
  wire [63:0] regs_424_io_out;
  wire  regs_424_io_enable;
  wire  regs_425_clock;
  wire  regs_425_reset;
  wire [63:0] regs_425_io_in;
  wire [63:0] regs_425_io_init;
  wire [63:0] regs_425_io_out;
  wire  regs_425_io_enable;
  wire  regs_426_clock;
  wire  regs_426_reset;
  wire [63:0] regs_426_io_in;
  wire [63:0] regs_426_io_init;
  wire [63:0] regs_426_io_out;
  wire  regs_426_io_enable;
  wire  regs_427_clock;
  wire  regs_427_reset;
  wire [63:0] regs_427_io_in;
  wire [63:0] regs_427_io_init;
  wire [63:0] regs_427_io_out;
  wire  regs_427_io_enable;
  wire  regs_428_clock;
  wire  regs_428_reset;
  wire [63:0] regs_428_io_in;
  wire [63:0] regs_428_io_init;
  wire [63:0] regs_428_io_out;
  wire  regs_428_io_enable;
  wire  regs_429_clock;
  wire  regs_429_reset;
  wire [63:0] regs_429_io_in;
  wire [63:0] regs_429_io_init;
  wire [63:0] regs_429_io_out;
  wire  regs_429_io_enable;
  wire  regs_430_clock;
  wire  regs_430_reset;
  wire [63:0] regs_430_io_in;
  wire [63:0] regs_430_io_init;
  wire [63:0] regs_430_io_out;
  wire  regs_430_io_enable;
  wire  regs_431_clock;
  wire  regs_431_reset;
  wire [63:0] regs_431_io_in;
  wire [63:0] regs_431_io_init;
  wire [63:0] regs_431_io_out;
  wire  regs_431_io_enable;
  wire  regs_432_clock;
  wire  regs_432_reset;
  wire [63:0] regs_432_io_in;
  wire [63:0] regs_432_io_init;
  wire [63:0] regs_432_io_out;
  wire  regs_432_io_enable;
  wire  regs_433_clock;
  wire  regs_433_reset;
  wire [63:0] regs_433_io_in;
  wire [63:0] regs_433_io_init;
  wire [63:0] regs_433_io_out;
  wire  regs_433_io_enable;
  wire  regs_434_clock;
  wire  regs_434_reset;
  wire [63:0] regs_434_io_in;
  wire [63:0] regs_434_io_init;
  wire [63:0] regs_434_io_out;
  wire  regs_434_io_enable;
  wire  regs_435_clock;
  wire  regs_435_reset;
  wire [63:0] regs_435_io_in;
  wire [63:0] regs_435_io_init;
  wire [63:0] regs_435_io_out;
  wire  regs_435_io_enable;
  wire  regs_436_clock;
  wire  regs_436_reset;
  wire [63:0] regs_436_io_in;
  wire [63:0] regs_436_io_init;
  wire [63:0] regs_436_io_out;
  wire  regs_436_io_enable;
  wire  regs_437_clock;
  wire  regs_437_reset;
  wire [63:0] regs_437_io_in;
  wire [63:0] regs_437_io_init;
  wire [63:0] regs_437_io_out;
  wire  regs_437_io_enable;
  wire  regs_438_clock;
  wire  regs_438_reset;
  wire [63:0] regs_438_io_in;
  wire [63:0] regs_438_io_init;
  wire [63:0] regs_438_io_out;
  wire  regs_438_io_enable;
  wire  regs_439_clock;
  wire  regs_439_reset;
  wire [63:0] regs_439_io_in;
  wire [63:0] regs_439_io_init;
  wire [63:0] regs_439_io_out;
  wire  regs_439_io_enable;
  wire  regs_440_clock;
  wire  regs_440_reset;
  wire [63:0] regs_440_io_in;
  wire [63:0] regs_440_io_init;
  wire [63:0] regs_440_io_out;
  wire  regs_440_io_enable;
  wire  regs_441_clock;
  wire  regs_441_reset;
  wire [63:0] regs_441_io_in;
  wire [63:0] regs_441_io_init;
  wire [63:0] regs_441_io_out;
  wire  regs_441_io_enable;
  wire  regs_442_clock;
  wire  regs_442_reset;
  wire [63:0] regs_442_io_in;
  wire [63:0] regs_442_io_init;
  wire [63:0] regs_442_io_out;
  wire  regs_442_io_enable;
  wire  regs_443_clock;
  wire  regs_443_reset;
  wire [63:0] regs_443_io_in;
  wire [63:0] regs_443_io_init;
  wire [63:0] regs_443_io_out;
  wire  regs_443_io_enable;
  wire  regs_444_clock;
  wire  regs_444_reset;
  wire [63:0] regs_444_io_in;
  wire [63:0] regs_444_io_init;
  wire [63:0] regs_444_io_out;
  wire  regs_444_io_enable;
  wire  regs_445_clock;
  wire  regs_445_reset;
  wire [63:0] regs_445_io_in;
  wire [63:0] regs_445_io_init;
  wire [63:0] regs_445_io_out;
  wire  regs_445_io_enable;
  wire  regs_446_clock;
  wire  regs_446_reset;
  wire [63:0] regs_446_io_in;
  wire [63:0] regs_446_io_init;
  wire [63:0] regs_446_io_out;
  wire  regs_446_io_enable;
  wire  regs_447_clock;
  wire  regs_447_reset;
  wire [63:0] regs_447_io_in;
  wire [63:0] regs_447_io_init;
  wire [63:0] regs_447_io_out;
  wire  regs_447_io_enable;
  wire  regs_448_clock;
  wire  regs_448_reset;
  wire [63:0] regs_448_io_in;
  wire [63:0] regs_448_io_init;
  wire [63:0] regs_448_io_out;
  wire  regs_448_io_enable;
  wire  regs_449_clock;
  wire  regs_449_reset;
  wire [63:0] regs_449_io_in;
  wire [63:0] regs_449_io_init;
  wire [63:0] regs_449_io_out;
  wire  regs_449_io_enable;
  wire  regs_450_clock;
  wire  regs_450_reset;
  wire [63:0] regs_450_io_in;
  wire [63:0] regs_450_io_init;
  wire [63:0] regs_450_io_out;
  wire  regs_450_io_enable;
  wire  regs_451_clock;
  wire  regs_451_reset;
  wire [63:0] regs_451_io_in;
  wire [63:0] regs_451_io_init;
  wire [63:0] regs_451_io_out;
  wire  regs_451_io_enable;
  wire  regs_452_clock;
  wire  regs_452_reset;
  wire [63:0] regs_452_io_in;
  wire [63:0] regs_452_io_init;
  wire [63:0] regs_452_io_out;
  wire  regs_452_io_enable;
  wire  regs_453_clock;
  wire  regs_453_reset;
  wire [63:0] regs_453_io_in;
  wire [63:0] regs_453_io_init;
  wire [63:0] regs_453_io_out;
  wire  regs_453_io_enable;
  wire  regs_454_clock;
  wire  regs_454_reset;
  wire [63:0] regs_454_io_in;
  wire [63:0] regs_454_io_init;
  wire [63:0] regs_454_io_out;
  wire  regs_454_io_enable;
  wire  regs_455_clock;
  wire  regs_455_reset;
  wire [63:0] regs_455_io_in;
  wire [63:0] regs_455_io_init;
  wire [63:0] regs_455_io_out;
  wire  regs_455_io_enable;
  wire  regs_456_clock;
  wire  regs_456_reset;
  wire [63:0] regs_456_io_in;
  wire [63:0] regs_456_io_init;
  wire [63:0] regs_456_io_out;
  wire  regs_456_io_enable;
  wire  regs_457_clock;
  wire  regs_457_reset;
  wire [63:0] regs_457_io_in;
  wire [63:0] regs_457_io_init;
  wire [63:0] regs_457_io_out;
  wire  regs_457_io_enable;
  wire  regs_458_clock;
  wire  regs_458_reset;
  wire [63:0] regs_458_io_in;
  wire [63:0] regs_458_io_init;
  wire [63:0] regs_458_io_out;
  wire  regs_458_io_enable;
  wire  regs_459_clock;
  wire  regs_459_reset;
  wire [63:0] regs_459_io_in;
  wire [63:0] regs_459_io_init;
  wire [63:0] regs_459_io_out;
  wire  regs_459_io_enable;
  wire  regs_460_clock;
  wire  regs_460_reset;
  wire [63:0] regs_460_io_in;
  wire [63:0] regs_460_io_init;
  wire [63:0] regs_460_io_out;
  wire  regs_460_io_enable;
  wire  regs_461_clock;
  wire  regs_461_reset;
  wire [63:0] regs_461_io_in;
  wire [63:0] regs_461_io_init;
  wire [63:0] regs_461_io_out;
  wire  regs_461_io_enable;
  wire  regs_462_clock;
  wire  regs_462_reset;
  wire [63:0] regs_462_io_in;
  wire [63:0] regs_462_io_init;
  wire [63:0] regs_462_io_out;
  wire  regs_462_io_enable;
  wire  regs_463_clock;
  wire  regs_463_reset;
  wire [63:0] regs_463_io_in;
  wire [63:0] regs_463_io_init;
  wire [63:0] regs_463_io_out;
  wire  regs_463_io_enable;
  wire  regs_464_clock;
  wire  regs_464_reset;
  wire [63:0] regs_464_io_in;
  wire [63:0] regs_464_io_init;
  wire [63:0] regs_464_io_out;
  wire  regs_464_io_enable;
  wire  regs_465_clock;
  wire  regs_465_reset;
  wire [63:0] regs_465_io_in;
  wire [63:0] regs_465_io_init;
  wire [63:0] regs_465_io_out;
  wire  regs_465_io_enable;
  wire  regs_466_clock;
  wire  regs_466_reset;
  wire [63:0] regs_466_io_in;
  wire [63:0] regs_466_io_init;
  wire [63:0] regs_466_io_out;
  wire  regs_466_io_enable;
  wire  regs_467_clock;
  wire  regs_467_reset;
  wire [63:0] regs_467_io_in;
  wire [63:0] regs_467_io_init;
  wire [63:0] regs_467_io_out;
  wire  regs_467_io_enable;
  wire  regs_468_clock;
  wire  regs_468_reset;
  wire [63:0] regs_468_io_in;
  wire [63:0] regs_468_io_init;
  wire [63:0] regs_468_io_out;
  wire  regs_468_io_enable;
  wire  regs_469_clock;
  wire  regs_469_reset;
  wire [63:0] regs_469_io_in;
  wire [63:0] regs_469_io_init;
  wire [63:0] regs_469_io_out;
  wire  regs_469_io_enable;
  wire  regs_470_clock;
  wire  regs_470_reset;
  wire [63:0] regs_470_io_in;
  wire [63:0] regs_470_io_init;
  wire [63:0] regs_470_io_out;
  wire  regs_470_io_enable;
  wire  regs_471_clock;
  wire  regs_471_reset;
  wire [63:0] regs_471_io_in;
  wire [63:0] regs_471_io_init;
  wire [63:0] regs_471_io_out;
  wire  regs_471_io_enable;
  wire  regs_472_clock;
  wire  regs_472_reset;
  wire [63:0] regs_472_io_in;
  wire [63:0] regs_472_io_init;
  wire [63:0] regs_472_io_out;
  wire  regs_472_io_enable;
  wire  regs_473_clock;
  wire  regs_473_reset;
  wire [63:0] regs_473_io_in;
  wire [63:0] regs_473_io_init;
  wire [63:0] regs_473_io_out;
  wire  regs_473_io_enable;
  wire  regs_474_clock;
  wire  regs_474_reset;
  wire [63:0] regs_474_io_in;
  wire [63:0] regs_474_io_init;
  wire [63:0] regs_474_io_out;
  wire  regs_474_io_enable;
  wire  regs_475_clock;
  wire  regs_475_reset;
  wire [63:0] regs_475_io_in;
  wire [63:0] regs_475_io_init;
  wire [63:0] regs_475_io_out;
  wire  regs_475_io_enable;
  wire  regs_476_clock;
  wire  regs_476_reset;
  wire [63:0] regs_476_io_in;
  wire [63:0] regs_476_io_init;
  wire [63:0] regs_476_io_out;
  wire  regs_476_io_enable;
  wire  regs_477_clock;
  wire  regs_477_reset;
  wire [63:0] regs_477_io_in;
  wire [63:0] regs_477_io_init;
  wire [63:0] regs_477_io_out;
  wire  regs_477_io_enable;
  wire  regs_478_clock;
  wire  regs_478_reset;
  wire [63:0] regs_478_io_in;
  wire [63:0] regs_478_io_init;
  wire [63:0] regs_478_io_out;
  wire  regs_478_io_enable;
  wire  regs_479_clock;
  wire  regs_479_reset;
  wire [63:0] regs_479_io_in;
  wire [63:0] regs_479_io_init;
  wire [63:0] regs_479_io_out;
  wire  regs_479_io_enable;
  wire  regs_480_clock;
  wire  regs_480_reset;
  wire [63:0] regs_480_io_in;
  wire [63:0] regs_480_io_init;
  wire [63:0] regs_480_io_out;
  wire  regs_480_io_enable;
  wire  regs_481_clock;
  wire  regs_481_reset;
  wire [63:0] regs_481_io_in;
  wire [63:0] regs_481_io_init;
  wire [63:0] regs_481_io_out;
  wire  regs_481_io_enable;
  wire  regs_482_clock;
  wire  regs_482_reset;
  wire [63:0] regs_482_io_in;
  wire [63:0] regs_482_io_init;
  wire [63:0] regs_482_io_out;
  wire  regs_482_io_enable;
  wire  regs_483_clock;
  wire  regs_483_reset;
  wire [63:0] regs_483_io_in;
  wire [63:0] regs_483_io_init;
  wire [63:0] regs_483_io_out;
  wire  regs_483_io_enable;
  wire  regs_484_clock;
  wire  regs_484_reset;
  wire [63:0] regs_484_io_in;
  wire [63:0] regs_484_io_init;
  wire [63:0] regs_484_io_out;
  wire  regs_484_io_enable;
  wire  regs_485_clock;
  wire  regs_485_reset;
  wire [63:0] regs_485_io_in;
  wire [63:0] regs_485_io_init;
  wire [63:0] regs_485_io_out;
  wire  regs_485_io_enable;
  wire  regs_486_clock;
  wire  regs_486_reset;
  wire [63:0] regs_486_io_in;
  wire [63:0] regs_486_io_init;
  wire [63:0] regs_486_io_out;
  wire  regs_486_io_enable;
  wire  regs_487_clock;
  wire  regs_487_reset;
  wire [63:0] regs_487_io_in;
  wire [63:0] regs_487_io_init;
  wire [63:0] regs_487_io_out;
  wire  regs_487_io_enable;
  wire  regs_488_clock;
  wire  regs_488_reset;
  wire [63:0] regs_488_io_in;
  wire [63:0] regs_488_io_init;
  wire [63:0] regs_488_io_out;
  wire  regs_488_io_enable;
  wire  regs_489_clock;
  wire  regs_489_reset;
  wire [63:0] regs_489_io_in;
  wire [63:0] regs_489_io_init;
  wire [63:0] regs_489_io_out;
  wire  regs_489_io_enable;
  wire  regs_490_clock;
  wire  regs_490_reset;
  wire [63:0] regs_490_io_in;
  wire [63:0] regs_490_io_init;
  wire [63:0] regs_490_io_out;
  wire  regs_490_io_enable;
  wire  regs_491_clock;
  wire  regs_491_reset;
  wire [63:0] regs_491_io_in;
  wire [63:0] regs_491_io_init;
  wire [63:0] regs_491_io_out;
  wire  regs_491_io_enable;
  wire  regs_492_clock;
  wire  regs_492_reset;
  wire [63:0] regs_492_io_in;
  wire [63:0] regs_492_io_init;
  wire [63:0] regs_492_io_out;
  wire  regs_492_io_enable;
  wire  regs_493_clock;
  wire  regs_493_reset;
  wire [63:0] regs_493_io_in;
  wire [63:0] regs_493_io_init;
  wire [63:0] regs_493_io_out;
  wire  regs_493_io_enable;
  wire  regs_494_clock;
  wire  regs_494_reset;
  wire [63:0] regs_494_io_in;
  wire [63:0] regs_494_io_init;
  wire [63:0] regs_494_io_out;
  wire  regs_494_io_enable;
  wire  regs_495_clock;
  wire  regs_495_reset;
  wire [63:0] regs_495_io_in;
  wire [63:0] regs_495_io_init;
  wire [63:0] regs_495_io_out;
  wire  regs_495_io_enable;
  wire  regs_496_clock;
  wire  regs_496_reset;
  wire [63:0] regs_496_io_in;
  wire [63:0] regs_496_io_init;
  wire [63:0] regs_496_io_out;
  wire  regs_496_io_enable;
  wire  regs_497_clock;
  wire  regs_497_reset;
  wire [63:0] regs_497_io_in;
  wire [63:0] regs_497_io_init;
  wire [63:0] regs_497_io_out;
  wire  regs_497_io_enable;
  wire  regs_498_clock;
  wire  regs_498_reset;
  wire [63:0] regs_498_io_in;
  wire [63:0] regs_498_io_init;
  wire [63:0] regs_498_io_out;
  wire  regs_498_io_enable;
  wire  regs_499_clock;
  wire  regs_499_reset;
  wire [63:0] regs_499_io_in;
  wire [63:0] regs_499_io_init;
  wire [63:0] regs_499_io_out;
  wire  regs_499_io_enable;
  wire  regs_500_clock;
  wire  regs_500_reset;
  wire [63:0] regs_500_io_in;
  wire [63:0] regs_500_io_init;
  wire [63:0] regs_500_io_out;
  wire  regs_500_io_enable;
  wire  regs_501_clock;
  wire  regs_501_reset;
  wire [63:0] regs_501_io_in;
  wire [63:0] regs_501_io_init;
  wire [63:0] regs_501_io_out;
  wire  regs_501_io_enable;
  wire  regs_502_clock;
  wire  regs_502_reset;
  wire [63:0] regs_502_io_in;
  wire [63:0] regs_502_io_init;
  wire [63:0] regs_502_io_out;
  wire  regs_502_io_enable;
  wire  regs_503_clock;
  wire  regs_503_reset;
  wire [63:0] regs_503_io_in;
  wire [63:0] regs_503_io_init;
  wire [63:0] regs_503_io_out;
  wire  regs_503_io_enable;
  wire  regs_504_clock;
  wire  regs_504_reset;
  wire [63:0] regs_504_io_in;
  wire [63:0] regs_504_io_init;
  wire [63:0] regs_504_io_out;
  wire  regs_504_io_enable;
  wire [63:0] rport_io_ins_0;
  wire [63:0] rport_io_ins_1;
  wire [63:0] rport_io_ins_2;
  wire [63:0] rport_io_ins_3;
  wire [63:0] rport_io_ins_4;
  wire [63:0] rport_io_ins_5;
  wire [63:0] rport_io_ins_6;
  wire [63:0] rport_io_ins_7;
  wire [63:0] rport_io_ins_8;
  wire [63:0] rport_io_ins_9;
  wire [63:0] rport_io_ins_10;
  wire [63:0] rport_io_ins_11;
  wire [63:0] rport_io_ins_12;
  wire [63:0] rport_io_ins_13;
  wire [63:0] rport_io_ins_14;
  wire [63:0] rport_io_ins_15;
  wire [63:0] rport_io_ins_16;
  wire [63:0] rport_io_ins_17;
  wire [63:0] rport_io_ins_18;
  wire [63:0] rport_io_ins_19;
  wire [63:0] rport_io_ins_20;
  wire [63:0] rport_io_ins_21;
  wire [63:0] rport_io_ins_22;
  wire [63:0] rport_io_ins_23;
  wire [63:0] rport_io_ins_24;
  wire [63:0] rport_io_ins_25;
  wire [63:0] rport_io_ins_26;
  wire [63:0] rport_io_ins_27;
  wire [63:0] rport_io_ins_28;
  wire [63:0] rport_io_ins_29;
  wire [63:0] rport_io_ins_30;
  wire [63:0] rport_io_ins_31;
  wire [63:0] rport_io_ins_32;
  wire [63:0] rport_io_ins_33;
  wire [63:0] rport_io_ins_34;
  wire [63:0] rport_io_ins_35;
  wire [63:0] rport_io_ins_36;
  wire [63:0] rport_io_ins_37;
  wire [63:0] rport_io_ins_38;
  wire [63:0] rport_io_ins_39;
  wire [63:0] rport_io_ins_40;
  wire [63:0] rport_io_ins_41;
  wire [63:0] rport_io_ins_42;
  wire [63:0] rport_io_ins_43;
  wire [63:0] rport_io_ins_44;
  wire [63:0] rport_io_ins_45;
  wire [63:0] rport_io_ins_46;
  wire [63:0] rport_io_ins_47;
  wire [63:0] rport_io_ins_48;
  wire [63:0] rport_io_ins_49;
  wire [63:0] rport_io_ins_50;
  wire [63:0] rport_io_ins_51;
  wire [63:0] rport_io_ins_52;
  wire [63:0] rport_io_ins_53;
  wire [63:0] rport_io_ins_54;
  wire [63:0] rport_io_ins_55;
  wire [63:0] rport_io_ins_56;
  wire [63:0] rport_io_ins_57;
  wire [63:0] rport_io_ins_58;
  wire [63:0] rport_io_ins_59;
  wire [63:0] rport_io_ins_60;
  wire [63:0] rport_io_ins_61;
  wire [63:0] rport_io_ins_62;
  wire [63:0] rport_io_ins_63;
  wire [63:0] rport_io_ins_64;
  wire [63:0] rport_io_ins_65;
  wire [63:0] rport_io_ins_66;
  wire [63:0] rport_io_ins_67;
  wire [63:0] rport_io_ins_68;
  wire [63:0] rport_io_ins_69;
  wire [63:0] rport_io_ins_70;
  wire [63:0] rport_io_ins_71;
  wire [63:0] rport_io_ins_72;
  wire [63:0] rport_io_ins_73;
  wire [63:0] rport_io_ins_74;
  wire [63:0] rport_io_ins_75;
  wire [63:0] rport_io_ins_76;
  wire [63:0] rport_io_ins_77;
  wire [63:0] rport_io_ins_78;
  wire [63:0] rport_io_ins_79;
  wire [63:0] rport_io_ins_80;
  wire [63:0] rport_io_ins_81;
  wire [63:0] rport_io_ins_82;
  wire [63:0] rport_io_ins_83;
  wire [63:0] rport_io_ins_84;
  wire [63:0] rport_io_ins_85;
  wire [63:0] rport_io_ins_86;
  wire [63:0] rport_io_ins_87;
  wire [63:0] rport_io_ins_88;
  wire [63:0] rport_io_ins_89;
  wire [63:0] rport_io_ins_90;
  wire [63:0] rport_io_ins_91;
  wire [63:0] rport_io_ins_92;
  wire [63:0] rport_io_ins_93;
  wire [63:0] rport_io_ins_94;
  wire [63:0] rport_io_ins_95;
  wire [63:0] rport_io_ins_96;
  wire [63:0] rport_io_ins_97;
  wire [63:0] rport_io_ins_98;
  wire [63:0] rport_io_ins_99;
  wire [63:0] rport_io_ins_100;
  wire [63:0] rport_io_ins_101;
  wire [63:0] rport_io_ins_102;
  wire [63:0] rport_io_ins_103;
  wire [63:0] rport_io_ins_104;
  wire [63:0] rport_io_ins_105;
  wire [63:0] rport_io_ins_106;
  wire [63:0] rport_io_ins_107;
  wire [63:0] rport_io_ins_108;
  wire [63:0] rport_io_ins_109;
  wire [63:0] rport_io_ins_110;
  wire [63:0] rport_io_ins_111;
  wire [63:0] rport_io_ins_112;
  wire [63:0] rport_io_ins_113;
  wire [63:0] rport_io_ins_114;
  wire [63:0] rport_io_ins_115;
  wire [63:0] rport_io_ins_116;
  wire [63:0] rport_io_ins_117;
  wire [63:0] rport_io_ins_118;
  wire [63:0] rport_io_ins_119;
  wire [63:0] rport_io_ins_120;
  wire [63:0] rport_io_ins_121;
  wire [63:0] rport_io_ins_122;
  wire [63:0] rport_io_ins_123;
  wire [63:0] rport_io_ins_124;
  wire [63:0] rport_io_ins_125;
  wire [63:0] rport_io_ins_126;
  wire [63:0] rport_io_ins_127;
  wire [63:0] rport_io_ins_128;
  wire [63:0] rport_io_ins_129;
  wire [63:0] rport_io_ins_130;
  wire [63:0] rport_io_ins_131;
  wire [63:0] rport_io_ins_132;
  wire [63:0] rport_io_ins_133;
  wire [63:0] rport_io_ins_134;
  wire [63:0] rport_io_ins_135;
  wire [63:0] rport_io_ins_136;
  wire [63:0] rport_io_ins_137;
  wire [63:0] rport_io_ins_138;
  wire [63:0] rport_io_ins_139;
  wire [63:0] rport_io_ins_140;
  wire [63:0] rport_io_ins_141;
  wire [63:0] rport_io_ins_142;
  wire [63:0] rport_io_ins_143;
  wire [63:0] rport_io_ins_144;
  wire [63:0] rport_io_ins_145;
  wire [63:0] rport_io_ins_146;
  wire [63:0] rport_io_ins_147;
  wire [63:0] rport_io_ins_148;
  wire [63:0] rport_io_ins_149;
  wire [63:0] rport_io_ins_150;
  wire [63:0] rport_io_ins_151;
  wire [63:0] rport_io_ins_152;
  wire [63:0] rport_io_ins_153;
  wire [63:0] rport_io_ins_154;
  wire [63:0] rport_io_ins_155;
  wire [63:0] rport_io_ins_156;
  wire [63:0] rport_io_ins_157;
  wire [63:0] rport_io_ins_158;
  wire [63:0] rport_io_ins_159;
  wire [63:0] rport_io_ins_160;
  wire [63:0] rport_io_ins_161;
  wire [63:0] rport_io_ins_162;
  wire [63:0] rport_io_ins_163;
  wire [63:0] rport_io_ins_164;
  wire [63:0] rport_io_ins_165;
  wire [63:0] rport_io_ins_166;
  wire [63:0] rport_io_ins_167;
  wire [63:0] rport_io_ins_168;
  wire [63:0] rport_io_ins_169;
  wire [63:0] rport_io_ins_170;
  wire [63:0] rport_io_ins_171;
  wire [63:0] rport_io_ins_172;
  wire [63:0] rport_io_ins_173;
  wire [63:0] rport_io_ins_174;
  wire [63:0] rport_io_ins_175;
  wire [63:0] rport_io_ins_176;
  wire [63:0] rport_io_ins_177;
  wire [63:0] rport_io_ins_178;
  wire [63:0] rport_io_ins_179;
  wire [63:0] rport_io_ins_180;
  wire [63:0] rport_io_ins_181;
  wire [63:0] rport_io_ins_182;
  wire [63:0] rport_io_ins_183;
  wire [63:0] rport_io_ins_184;
  wire [63:0] rport_io_ins_185;
  wire [63:0] rport_io_ins_186;
  wire [63:0] rport_io_ins_187;
  wire [63:0] rport_io_ins_188;
  wire [63:0] rport_io_ins_189;
  wire [63:0] rport_io_ins_190;
  wire [63:0] rport_io_ins_191;
  wire [63:0] rport_io_ins_192;
  wire [63:0] rport_io_ins_193;
  wire [63:0] rport_io_ins_194;
  wire [63:0] rport_io_ins_195;
  wire [63:0] rport_io_ins_196;
  wire [63:0] rport_io_ins_197;
  wire [63:0] rport_io_ins_198;
  wire [63:0] rport_io_ins_199;
  wire [63:0] rport_io_ins_200;
  wire [63:0] rport_io_ins_201;
  wire [63:0] rport_io_ins_202;
  wire [63:0] rport_io_ins_203;
  wire [63:0] rport_io_ins_204;
  wire [63:0] rport_io_ins_205;
  wire [63:0] rport_io_ins_206;
  wire [63:0] rport_io_ins_207;
  wire [63:0] rport_io_ins_208;
  wire [63:0] rport_io_ins_209;
  wire [63:0] rport_io_ins_210;
  wire [63:0] rport_io_ins_211;
  wire [63:0] rport_io_ins_212;
  wire [63:0] rport_io_ins_213;
  wire [63:0] rport_io_ins_214;
  wire [63:0] rport_io_ins_215;
  wire [63:0] rport_io_ins_216;
  wire [63:0] rport_io_ins_217;
  wire [63:0] rport_io_ins_218;
  wire [63:0] rport_io_ins_219;
  wire [63:0] rport_io_ins_220;
  wire [63:0] rport_io_ins_221;
  wire [63:0] rport_io_ins_222;
  wire [63:0] rport_io_ins_223;
  wire [63:0] rport_io_ins_224;
  wire [63:0] rport_io_ins_225;
  wire [63:0] rport_io_ins_226;
  wire [63:0] rport_io_ins_227;
  wire [63:0] rport_io_ins_228;
  wire [63:0] rport_io_ins_229;
  wire [63:0] rport_io_ins_230;
  wire [63:0] rport_io_ins_231;
  wire [63:0] rport_io_ins_232;
  wire [63:0] rport_io_ins_233;
  wire [63:0] rport_io_ins_234;
  wire [63:0] rport_io_ins_235;
  wire [63:0] rport_io_ins_236;
  wire [63:0] rport_io_ins_237;
  wire [63:0] rport_io_ins_238;
  wire [63:0] rport_io_ins_239;
  wire [63:0] rport_io_ins_240;
  wire [63:0] rport_io_ins_241;
  wire [63:0] rport_io_ins_242;
  wire [63:0] rport_io_ins_243;
  wire [63:0] rport_io_ins_244;
  wire [63:0] rport_io_ins_245;
  wire [63:0] rport_io_ins_246;
  wire [63:0] rport_io_ins_247;
  wire [63:0] rport_io_ins_248;
  wire [63:0] rport_io_ins_249;
  wire [63:0] rport_io_ins_250;
  wire [63:0] rport_io_ins_251;
  wire [63:0] rport_io_ins_252;
  wire [63:0] rport_io_ins_253;
  wire [63:0] rport_io_ins_254;
  wire [63:0] rport_io_ins_255;
  wire [63:0] rport_io_ins_256;
  wire [63:0] rport_io_ins_257;
  wire [63:0] rport_io_ins_258;
  wire [63:0] rport_io_ins_259;
  wire [63:0] rport_io_ins_260;
  wire [63:0] rport_io_ins_261;
  wire [63:0] rport_io_ins_262;
  wire [63:0] rport_io_ins_263;
  wire [63:0] rport_io_ins_264;
  wire [63:0] rport_io_ins_265;
  wire [63:0] rport_io_ins_266;
  wire [63:0] rport_io_ins_267;
  wire [63:0] rport_io_ins_268;
  wire [63:0] rport_io_ins_269;
  wire [63:0] rport_io_ins_270;
  wire [63:0] rport_io_ins_271;
  wire [63:0] rport_io_ins_272;
  wire [63:0] rport_io_ins_273;
  wire [63:0] rport_io_ins_274;
  wire [63:0] rport_io_ins_275;
  wire [63:0] rport_io_ins_276;
  wire [63:0] rport_io_ins_277;
  wire [63:0] rport_io_ins_278;
  wire [63:0] rport_io_ins_279;
  wire [63:0] rport_io_ins_280;
  wire [63:0] rport_io_ins_281;
  wire [63:0] rport_io_ins_282;
  wire [63:0] rport_io_ins_283;
  wire [63:0] rport_io_ins_284;
  wire [63:0] rport_io_ins_285;
  wire [63:0] rport_io_ins_286;
  wire [63:0] rport_io_ins_287;
  wire [63:0] rport_io_ins_288;
  wire [63:0] rport_io_ins_289;
  wire [63:0] rport_io_ins_290;
  wire [63:0] rport_io_ins_291;
  wire [63:0] rport_io_ins_292;
  wire [63:0] rport_io_ins_293;
  wire [63:0] rport_io_ins_294;
  wire [63:0] rport_io_ins_295;
  wire [63:0] rport_io_ins_296;
  wire [63:0] rport_io_ins_297;
  wire [63:0] rport_io_ins_298;
  wire [63:0] rport_io_ins_299;
  wire [63:0] rport_io_ins_300;
  wire [63:0] rport_io_ins_301;
  wire [63:0] rport_io_ins_302;
  wire [63:0] rport_io_ins_303;
  wire [63:0] rport_io_ins_304;
  wire [63:0] rport_io_ins_305;
  wire [63:0] rport_io_ins_306;
  wire [63:0] rport_io_ins_307;
  wire [63:0] rport_io_ins_308;
  wire [63:0] rport_io_ins_309;
  wire [63:0] rport_io_ins_310;
  wire [63:0] rport_io_ins_311;
  wire [63:0] rport_io_ins_312;
  wire [63:0] rport_io_ins_313;
  wire [63:0] rport_io_ins_314;
  wire [63:0] rport_io_ins_315;
  wire [63:0] rport_io_ins_316;
  wire [63:0] rport_io_ins_317;
  wire [63:0] rport_io_ins_318;
  wire [63:0] rport_io_ins_319;
  wire [63:0] rport_io_ins_320;
  wire [63:0] rport_io_ins_321;
  wire [63:0] rport_io_ins_322;
  wire [63:0] rport_io_ins_323;
  wire [63:0] rport_io_ins_324;
  wire [63:0] rport_io_ins_325;
  wire [63:0] rport_io_ins_326;
  wire [63:0] rport_io_ins_327;
  wire [63:0] rport_io_ins_328;
  wire [63:0] rport_io_ins_329;
  wire [63:0] rport_io_ins_330;
  wire [63:0] rport_io_ins_331;
  wire [63:0] rport_io_ins_332;
  wire [63:0] rport_io_ins_333;
  wire [63:0] rport_io_ins_334;
  wire [63:0] rport_io_ins_335;
  wire [63:0] rport_io_ins_336;
  wire [63:0] rport_io_ins_337;
  wire [63:0] rport_io_ins_338;
  wire [63:0] rport_io_ins_339;
  wire [63:0] rport_io_ins_340;
  wire [63:0] rport_io_ins_341;
  wire [63:0] rport_io_ins_342;
  wire [63:0] rport_io_ins_343;
  wire [63:0] rport_io_ins_344;
  wire [63:0] rport_io_ins_345;
  wire [63:0] rport_io_ins_346;
  wire [63:0] rport_io_ins_347;
  wire [63:0] rport_io_ins_348;
  wire [63:0] rport_io_ins_349;
  wire [63:0] rport_io_ins_350;
  wire [63:0] rport_io_ins_351;
  wire [63:0] rport_io_ins_352;
  wire [63:0] rport_io_ins_353;
  wire [63:0] rport_io_ins_354;
  wire [63:0] rport_io_ins_355;
  wire [63:0] rport_io_ins_356;
  wire [63:0] rport_io_ins_357;
  wire [63:0] rport_io_ins_358;
  wire [63:0] rport_io_ins_359;
  wire [63:0] rport_io_ins_360;
  wire [63:0] rport_io_ins_361;
  wire [63:0] rport_io_ins_362;
  wire [63:0] rport_io_ins_363;
  wire [63:0] rport_io_ins_364;
  wire [63:0] rport_io_ins_365;
  wire [63:0] rport_io_ins_366;
  wire [63:0] rport_io_ins_367;
  wire [63:0] rport_io_ins_368;
  wire [63:0] rport_io_ins_369;
  wire [63:0] rport_io_ins_370;
  wire [63:0] rport_io_ins_371;
  wire [63:0] rport_io_ins_372;
  wire [63:0] rport_io_ins_373;
  wire [63:0] rport_io_ins_374;
  wire [63:0] rport_io_ins_375;
  wire [63:0] rport_io_ins_376;
  wire [63:0] rport_io_ins_377;
  wire [63:0] rport_io_ins_378;
  wire [63:0] rport_io_ins_379;
  wire [63:0] rport_io_ins_380;
  wire [63:0] rport_io_ins_381;
  wire [63:0] rport_io_ins_382;
  wire [63:0] rport_io_ins_383;
  wire [63:0] rport_io_ins_384;
  wire [63:0] rport_io_ins_385;
  wire [63:0] rport_io_ins_386;
  wire [63:0] rport_io_ins_387;
  wire [63:0] rport_io_ins_388;
  wire [63:0] rport_io_ins_389;
  wire [63:0] rport_io_ins_390;
  wire [63:0] rport_io_ins_391;
  wire [63:0] rport_io_ins_392;
  wire [63:0] rport_io_ins_393;
  wire [63:0] rport_io_ins_394;
  wire [63:0] rport_io_ins_395;
  wire [63:0] rport_io_ins_396;
  wire [63:0] rport_io_ins_397;
  wire [63:0] rport_io_ins_398;
  wire [63:0] rport_io_ins_399;
  wire [63:0] rport_io_ins_400;
  wire [63:0] rport_io_ins_401;
  wire [63:0] rport_io_ins_402;
  wire [63:0] rport_io_ins_403;
  wire [63:0] rport_io_ins_404;
  wire [63:0] rport_io_ins_405;
  wire [63:0] rport_io_ins_406;
  wire [63:0] rport_io_ins_407;
  wire [63:0] rport_io_ins_408;
  wire [63:0] rport_io_ins_409;
  wire [63:0] rport_io_ins_410;
  wire [63:0] rport_io_ins_411;
  wire [63:0] rport_io_ins_412;
  wire [63:0] rport_io_ins_413;
  wire [63:0] rport_io_ins_414;
  wire [63:0] rport_io_ins_415;
  wire [63:0] rport_io_ins_416;
  wire [63:0] rport_io_ins_417;
  wire [63:0] rport_io_ins_418;
  wire [63:0] rport_io_ins_419;
  wire [63:0] rport_io_ins_420;
  wire [63:0] rport_io_ins_421;
  wire [63:0] rport_io_ins_422;
  wire [63:0] rport_io_ins_423;
  wire [63:0] rport_io_ins_424;
  wire [63:0] rport_io_ins_425;
  wire [63:0] rport_io_ins_426;
  wire [63:0] rport_io_ins_427;
  wire [63:0] rport_io_ins_428;
  wire [63:0] rport_io_ins_429;
  wire [63:0] rport_io_ins_430;
  wire [63:0] rport_io_ins_431;
  wire [63:0] rport_io_ins_432;
  wire [63:0] rport_io_ins_433;
  wire [63:0] rport_io_ins_434;
  wire [63:0] rport_io_ins_435;
  wire [63:0] rport_io_ins_436;
  wire [63:0] rport_io_ins_437;
  wire [63:0] rport_io_ins_438;
  wire [63:0] rport_io_ins_439;
  wire [63:0] rport_io_ins_440;
  wire [63:0] rport_io_ins_441;
  wire [63:0] rport_io_ins_442;
  wire [63:0] rport_io_ins_443;
  wire [63:0] rport_io_ins_444;
  wire [63:0] rport_io_ins_445;
  wire [63:0] rport_io_ins_446;
  wire [63:0] rport_io_ins_447;
  wire [63:0] rport_io_ins_448;
  wire [63:0] rport_io_ins_449;
  wire [63:0] rport_io_ins_450;
  wire [63:0] rport_io_ins_451;
  wire [63:0] rport_io_ins_452;
  wire [63:0] rport_io_ins_453;
  wire [63:0] rport_io_ins_454;
  wire [63:0] rport_io_ins_455;
  wire [63:0] rport_io_ins_456;
  wire [63:0] rport_io_ins_457;
  wire [63:0] rport_io_ins_458;
  wire [63:0] rport_io_ins_459;
  wire [63:0] rport_io_ins_460;
  wire [63:0] rport_io_ins_461;
  wire [63:0] rport_io_ins_462;
  wire [63:0] rport_io_ins_463;
  wire [63:0] rport_io_ins_464;
  wire [63:0] rport_io_ins_465;
  wire [63:0] rport_io_ins_466;
  wire [63:0] rport_io_ins_467;
  wire [63:0] rport_io_ins_468;
  wire [63:0] rport_io_ins_469;
  wire [63:0] rport_io_ins_470;
  wire [63:0] rport_io_ins_471;
  wire [63:0] rport_io_ins_472;
  wire [63:0] rport_io_ins_473;
  wire [63:0] rport_io_ins_474;
  wire [63:0] rport_io_ins_475;
  wire [63:0] rport_io_ins_476;
  wire [63:0] rport_io_ins_477;
  wire [63:0] rport_io_ins_478;
  wire [63:0] rport_io_ins_479;
  wire [63:0] rport_io_ins_480;
  wire [63:0] rport_io_ins_481;
  wire [63:0] rport_io_ins_482;
  wire [63:0] rport_io_ins_483;
  wire [63:0] rport_io_ins_484;
  wire [63:0] rport_io_ins_485;
  wire [63:0] rport_io_ins_486;
  wire [63:0] rport_io_ins_487;
  wire [63:0] rport_io_ins_488;
  wire [63:0] rport_io_ins_489;
  wire [63:0] rport_io_ins_490;
  wire [63:0] rport_io_ins_491;
  wire [63:0] rport_io_ins_492;
  wire [63:0] rport_io_ins_493;
  wire [63:0] rport_io_ins_494;
  wire [63:0] rport_io_ins_495;
  wire [63:0] rport_io_ins_496;
  wire [63:0] rport_io_ins_497;
  wire [63:0] rport_io_ins_498;
  wire [63:0] rport_io_ins_499;
  wire [63:0] rport_io_ins_500;
  wire [63:0] rport_io_ins_501;
  wire [63:0] rport_io_ins_502;
  wire [63:0] rport_io_ins_503;
  wire [63:0] rport_io_ins_504;
  wire [8:0] rport_io_sel;
  wire [63:0] rport_io_out;
  wire [63:0] regOuts_0;
  wire [63:0] regOuts_1;
  wire [63:0] regOuts_2;
  wire [63:0] regOuts_3;
  wire [63:0] regOuts_4;
  wire [63:0] regOuts_5;
  wire [63:0] regOuts_6;
  wire [63:0] regOuts_7;
  wire [63:0] regOuts_8;
  wire [63:0] regOuts_9;
  wire [63:0] regOuts_10;
  wire [63:0] regOuts_11;
  wire [63:0] regOuts_12;
  wire [63:0] regOuts_13;
  wire [63:0] regOuts_14;
  wire [63:0] regOuts_15;
  wire [63:0] regOuts_16;
  wire [63:0] regOuts_17;
  wire [63:0] regOuts_18;
  wire [63:0] regOuts_19;
  wire [63:0] regOuts_20;
  wire [63:0] regOuts_21;
  wire [63:0] regOuts_22;
  wire [63:0] regOuts_23;
  wire [63:0] regOuts_24;
  wire [63:0] regOuts_25;
  wire [63:0] regOuts_26;
  wire [63:0] regOuts_27;
  wire [63:0] regOuts_28;
  wire [63:0] regOuts_29;
  wire [63:0] regOuts_30;
  wire [63:0] regOuts_31;
  wire [63:0] regOuts_32;
  wire [63:0] regOuts_33;
  wire [63:0] regOuts_34;
  wire [63:0] regOuts_35;
  wire [63:0] regOuts_36;
  wire [63:0] regOuts_37;
  wire [63:0] regOuts_38;
  wire [63:0] regOuts_39;
  wire [63:0] regOuts_40;
  wire [63:0] regOuts_41;
  wire [63:0] regOuts_42;
  wire [63:0] regOuts_43;
  wire [63:0] regOuts_44;
  wire [63:0] regOuts_45;
  wire [63:0] regOuts_46;
  wire [63:0] regOuts_47;
  wire [63:0] regOuts_48;
  wire [63:0] regOuts_49;
  wire [63:0] regOuts_50;
  wire [63:0] regOuts_51;
  wire [63:0] regOuts_52;
  wire [63:0] regOuts_53;
  wire [63:0] regOuts_54;
  wire [63:0] regOuts_55;
  wire [63:0] regOuts_56;
  wire [63:0] regOuts_57;
  wire [63:0] regOuts_58;
  wire [63:0] regOuts_59;
  wire [63:0] regOuts_60;
  wire [63:0] regOuts_61;
  wire [63:0] regOuts_62;
  wire [63:0] regOuts_63;
  wire [63:0] regOuts_64;
  wire [63:0] regOuts_65;
  wire [63:0] regOuts_66;
  wire [63:0] regOuts_67;
  wire [63:0] regOuts_68;
  wire [63:0] regOuts_69;
  wire [63:0] regOuts_70;
  wire [63:0] regOuts_71;
  wire [63:0] regOuts_72;
  wire [63:0] regOuts_73;
  wire [63:0] regOuts_74;
  wire [63:0] regOuts_75;
  wire [63:0] regOuts_76;
  wire [63:0] regOuts_77;
  wire [63:0] regOuts_78;
  wire [63:0] regOuts_79;
  wire [63:0] regOuts_80;
  wire [63:0] regOuts_81;
  wire [63:0] regOuts_82;
  wire [63:0] regOuts_83;
  wire [63:0] regOuts_84;
  wire [63:0] regOuts_85;
  wire [63:0] regOuts_86;
  wire [63:0] regOuts_87;
  wire [63:0] regOuts_88;
  wire [63:0] regOuts_89;
  wire [63:0] regOuts_90;
  wire [63:0] regOuts_91;
  wire [63:0] regOuts_92;
  wire [63:0] regOuts_93;
  wire [63:0] regOuts_94;
  wire [63:0] regOuts_95;
  wire [63:0] regOuts_96;
  wire [63:0] regOuts_97;
  wire [63:0] regOuts_98;
  wire [63:0] regOuts_99;
  wire [63:0] regOuts_100;
  wire [63:0] regOuts_101;
  wire [63:0] regOuts_102;
  wire [63:0] regOuts_103;
  wire [63:0] regOuts_104;
  wire [63:0] regOuts_105;
  wire [63:0] regOuts_106;
  wire [63:0] regOuts_107;
  wire [63:0] regOuts_108;
  wire [63:0] regOuts_109;
  wire [63:0] regOuts_110;
  wire [63:0] regOuts_111;
  wire [63:0] regOuts_112;
  wire [63:0] regOuts_113;
  wire [63:0] regOuts_114;
  wire [63:0] regOuts_115;
  wire [63:0] regOuts_116;
  wire [63:0] regOuts_117;
  wire [63:0] regOuts_118;
  wire [63:0] regOuts_119;
  wire [63:0] regOuts_120;
  wire [63:0] regOuts_121;
  wire [63:0] regOuts_122;
  wire [63:0] regOuts_123;
  wire [63:0] regOuts_124;
  wire [63:0] regOuts_125;
  wire [63:0] regOuts_126;
  wire [63:0] regOuts_127;
  wire [63:0] regOuts_128;
  wire [63:0] regOuts_129;
  wire [63:0] regOuts_130;
  wire [63:0] regOuts_131;
  wire [63:0] regOuts_132;
  wire [63:0] regOuts_133;
  wire [63:0] regOuts_134;
  wire [63:0] regOuts_135;
  wire [63:0] regOuts_136;
  wire [63:0] regOuts_137;
  wire [63:0] regOuts_138;
  wire [63:0] regOuts_139;
  wire [63:0] regOuts_140;
  wire [63:0] regOuts_141;
  wire [63:0] regOuts_142;
  wire [63:0] regOuts_143;
  wire [63:0] regOuts_144;
  wire [63:0] regOuts_145;
  wire [63:0] regOuts_146;
  wire [63:0] regOuts_147;
  wire [63:0] regOuts_148;
  wire [63:0] regOuts_149;
  wire [63:0] regOuts_150;
  wire [63:0] regOuts_151;
  wire [63:0] regOuts_152;
  wire [63:0] regOuts_153;
  wire [63:0] regOuts_154;
  wire [63:0] regOuts_155;
  wire [63:0] regOuts_156;
  wire [63:0] regOuts_157;
  wire [63:0] regOuts_158;
  wire [63:0] regOuts_159;
  wire [63:0] regOuts_160;
  wire [63:0] regOuts_161;
  wire [63:0] regOuts_162;
  wire [63:0] regOuts_163;
  wire [63:0] regOuts_164;
  wire [63:0] regOuts_165;
  wire [63:0] regOuts_166;
  wire [63:0] regOuts_167;
  wire [63:0] regOuts_168;
  wire [63:0] regOuts_169;
  wire [63:0] regOuts_170;
  wire [63:0] regOuts_171;
  wire [63:0] regOuts_172;
  wire [63:0] regOuts_173;
  wire [63:0] regOuts_174;
  wire [63:0] regOuts_175;
  wire [63:0] regOuts_176;
  wire [63:0] regOuts_177;
  wire [63:0] regOuts_178;
  wire [63:0] regOuts_179;
  wire [63:0] regOuts_180;
  wire [63:0] regOuts_181;
  wire [63:0] regOuts_182;
  wire [63:0] regOuts_183;
  wire [63:0] regOuts_184;
  wire [63:0] regOuts_185;
  wire [63:0] regOuts_186;
  wire [63:0] regOuts_187;
  wire [63:0] regOuts_188;
  wire [63:0] regOuts_189;
  wire [63:0] regOuts_190;
  wire [63:0] regOuts_191;
  wire [63:0] regOuts_192;
  wire [63:0] regOuts_193;
  wire [63:0] regOuts_194;
  wire [63:0] regOuts_195;
  wire [63:0] regOuts_196;
  wire [63:0] regOuts_197;
  wire [63:0] regOuts_198;
  wire [63:0] regOuts_199;
  wire [63:0] regOuts_200;
  wire [63:0] regOuts_201;
  wire [63:0] regOuts_202;
  wire [63:0] regOuts_203;
  wire [63:0] regOuts_204;
  wire [63:0] regOuts_205;
  wire [63:0] regOuts_206;
  wire [63:0] regOuts_207;
  wire [63:0] regOuts_208;
  wire [63:0] regOuts_209;
  wire [63:0] regOuts_210;
  wire [63:0] regOuts_211;
  wire [63:0] regOuts_212;
  wire [63:0] regOuts_213;
  wire [63:0] regOuts_214;
  wire [63:0] regOuts_215;
  wire [63:0] regOuts_216;
  wire [63:0] regOuts_217;
  wire [63:0] regOuts_218;
  wire [63:0] regOuts_219;
  wire [63:0] regOuts_220;
  wire [63:0] regOuts_221;
  wire [63:0] regOuts_222;
  wire [63:0] regOuts_223;
  wire [63:0] regOuts_224;
  wire [63:0] regOuts_225;
  wire [63:0] regOuts_226;
  wire [63:0] regOuts_227;
  wire [63:0] regOuts_228;
  wire [63:0] regOuts_229;
  wire [63:0] regOuts_230;
  wire [63:0] regOuts_231;
  wire [63:0] regOuts_232;
  wire [63:0] regOuts_233;
  wire [63:0] regOuts_234;
  wire [63:0] regOuts_235;
  wire [63:0] regOuts_236;
  wire [63:0] regOuts_237;
  wire [63:0] regOuts_238;
  wire [63:0] regOuts_239;
  wire [63:0] regOuts_240;
  wire [63:0] regOuts_241;
  wire [63:0] regOuts_242;
  wire [63:0] regOuts_243;
  wire [63:0] regOuts_244;
  wire [63:0] regOuts_245;
  wire [63:0] regOuts_246;
  wire [63:0] regOuts_247;
  wire [63:0] regOuts_248;
  wire [63:0] regOuts_249;
  wire [63:0] regOuts_250;
  wire [63:0] regOuts_251;
  wire [63:0] regOuts_252;
  wire [63:0] regOuts_253;
  wire [63:0] regOuts_254;
  wire [63:0] regOuts_255;
  wire [63:0] regOuts_256;
  wire [63:0] regOuts_257;
  wire [63:0] regOuts_258;
  wire [63:0] regOuts_259;
  wire [63:0] regOuts_260;
  wire [63:0] regOuts_261;
  wire [63:0] regOuts_262;
  wire [63:0] regOuts_263;
  wire [63:0] regOuts_264;
  wire [63:0] regOuts_265;
  wire [63:0] regOuts_266;
  wire [63:0] regOuts_267;
  wire [63:0] regOuts_268;
  wire [63:0] regOuts_269;
  wire [63:0] regOuts_270;
  wire [63:0] regOuts_271;
  wire [63:0] regOuts_272;
  wire [63:0] regOuts_273;
  wire [63:0] regOuts_274;
  wire [63:0] regOuts_275;
  wire [63:0] regOuts_276;
  wire [63:0] regOuts_277;
  wire [63:0] regOuts_278;
  wire [63:0] regOuts_279;
  wire [63:0] regOuts_280;
  wire [63:0] regOuts_281;
  wire [63:0] regOuts_282;
  wire [63:0] regOuts_283;
  wire [63:0] regOuts_284;
  wire [63:0] regOuts_285;
  wire [63:0] regOuts_286;
  wire [63:0] regOuts_287;
  wire [63:0] regOuts_288;
  wire [63:0] regOuts_289;
  wire [63:0] regOuts_290;
  wire [63:0] regOuts_291;
  wire [63:0] regOuts_292;
  wire [63:0] regOuts_293;
  wire [63:0] regOuts_294;
  wire [63:0] regOuts_295;
  wire [63:0] regOuts_296;
  wire [63:0] regOuts_297;
  wire [63:0] regOuts_298;
  wire [63:0] regOuts_299;
  wire [63:0] regOuts_300;
  wire [63:0] regOuts_301;
  wire [63:0] regOuts_302;
  wire [63:0] regOuts_303;
  wire [63:0] regOuts_304;
  wire [63:0] regOuts_305;
  wire [63:0] regOuts_306;
  wire [63:0] regOuts_307;
  wire [63:0] regOuts_308;
  wire [63:0] regOuts_309;
  wire [63:0] regOuts_310;
  wire [63:0] regOuts_311;
  wire [63:0] regOuts_312;
  wire [63:0] regOuts_313;
  wire [63:0] regOuts_314;
  wire [63:0] regOuts_315;
  wire [63:0] regOuts_316;
  wire [63:0] regOuts_317;
  wire [63:0] regOuts_318;
  wire [63:0] regOuts_319;
  wire [63:0] regOuts_320;
  wire [63:0] regOuts_321;
  wire [63:0] regOuts_322;
  wire [63:0] regOuts_323;
  wire [63:0] regOuts_324;
  wire [63:0] regOuts_325;
  wire [63:0] regOuts_326;
  wire [63:0] regOuts_327;
  wire [63:0] regOuts_328;
  wire [63:0] regOuts_329;
  wire [63:0] regOuts_330;
  wire [63:0] regOuts_331;
  wire [63:0] regOuts_332;
  wire [63:0] regOuts_333;
  wire [63:0] regOuts_334;
  wire [63:0] regOuts_335;
  wire [63:0] regOuts_336;
  wire [63:0] regOuts_337;
  wire [63:0] regOuts_338;
  wire [63:0] regOuts_339;
  wire [63:0] regOuts_340;
  wire [63:0] regOuts_341;
  wire [63:0] regOuts_342;
  wire [63:0] regOuts_343;
  wire [63:0] regOuts_344;
  wire [63:0] regOuts_345;
  wire [63:0] regOuts_346;
  wire [63:0] regOuts_347;
  wire [63:0] regOuts_348;
  wire [63:0] regOuts_349;
  wire [63:0] regOuts_350;
  wire [63:0] regOuts_351;
  wire [63:0] regOuts_352;
  wire [63:0] regOuts_353;
  wire [63:0] regOuts_354;
  wire [63:0] regOuts_355;
  wire [63:0] regOuts_356;
  wire [63:0] regOuts_357;
  wire [63:0] regOuts_358;
  wire [63:0] regOuts_359;
  wire [63:0] regOuts_360;
  wire [63:0] regOuts_361;
  wire [63:0] regOuts_362;
  wire [63:0] regOuts_363;
  wire [63:0] regOuts_364;
  wire [63:0] regOuts_365;
  wire [63:0] regOuts_366;
  wire [63:0] regOuts_367;
  wire [63:0] regOuts_368;
  wire [63:0] regOuts_369;
  wire [63:0] regOuts_370;
  wire [63:0] regOuts_371;
  wire [63:0] regOuts_372;
  wire [63:0] regOuts_373;
  wire [63:0] regOuts_374;
  wire [63:0] regOuts_375;
  wire [63:0] regOuts_376;
  wire [63:0] regOuts_377;
  wire [63:0] regOuts_378;
  wire [63:0] regOuts_379;
  wire [63:0] regOuts_380;
  wire [63:0] regOuts_381;
  wire [63:0] regOuts_382;
  wire [63:0] regOuts_383;
  wire [63:0] regOuts_384;
  wire [63:0] regOuts_385;
  wire [63:0] regOuts_386;
  wire [63:0] regOuts_387;
  wire [63:0] regOuts_388;
  wire [63:0] regOuts_389;
  wire [63:0] regOuts_390;
  wire [63:0] regOuts_391;
  wire [63:0] regOuts_392;
  wire [63:0] regOuts_393;
  wire [63:0] regOuts_394;
  wire [63:0] regOuts_395;
  wire [63:0] regOuts_396;
  wire [63:0] regOuts_397;
  wire [63:0] regOuts_398;
  wire [63:0] regOuts_399;
  wire [63:0] regOuts_400;
  wire [63:0] regOuts_401;
  wire [63:0] regOuts_402;
  wire [63:0] regOuts_403;
  wire [63:0] regOuts_404;
  wire [63:0] regOuts_405;
  wire [63:0] regOuts_406;
  wire [63:0] regOuts_407;
  wire [63:0] regOuts_408;
  wire [63:0] regOuts_409;
  wire [63:0] regOuts_410;
  wire [63:0] regOuts_411;
  wire [63:0] regOuts_412;
  wire [63:0] regOuts_413;
  wire [63:0] regOuts_414;
  wire [63:0] regOuts_415;
  wire [63:0] regOuts_416;
  wire [63:0] regOuts_417;
  wire [63:0] regOuts_418;
  wire [63:0] regOuts_419;
  wire [63:0] regOuts_420;
  wire [63:0] regOuts_421;
  wire [63:0] regOuts_422;
  wire [63:0] regOuts_423;
  wire [63:0] regOuts_424;
  wire [63:0] regOuts_425;
  wire [63:0] regOuts_426;
  wire [63:0] regOuts_427;
  wire [63:0] regOuts_428;
  wire [63:0] regOuts_429;
  wire [63:0] regOuts_430;
  wire [63:0] regOuts_431;
  wire [63:0] regOuts_432;
  wire [63:0] regOuts_433;
  wire [63:0] regOuts_434;
  wire [63:0] regOuts_435;
  wire [63:0] regOuts_436;
  wire [63:0] regOuts_437;
  wire [63:0] regOuts_438;
  wire [63:0] regOuts_439;
  wire [63:0] regOuts_440;
  wire [63:0] regOuts_441;
  wire [63:0] regOuts_442;
  wire [63:0] regOuts_443;
  wire [63:0] regOuts_444;
  wire [63:0] regOuts_445;
  wire [63:0] regOuts_446;
  wire [63:0] regOuts_447;
  wire [63:0] regOuts_448;
  wire [63:0] regOuts_449;
  wire [63:0] regOuts_450;
  wire [63:0] regOuts_451;
  wire [63:0] regOuts_452;
  wire [63:0] regOuts_453;
  wire [63:0] regOuts_454;
  wire [63:0] regOuts_455;
  wire [63:0] regOuts_456;
  wire [63:0] regOuts_457;
  wire [63:0] regOuts_458;
  wire [63:0] regOuts_459;
  wire [63:0] regOuts_460;
  wire [63:0] regOuts_461;
  wire [63:0] regOuts_462;
  wire [63:0] regOuts_463;
  wire [63:0] regOuts_464;
  wire [63:0] regOuts_465;
  wire [63:0] regOuts_466;
  wire [63:0] regOuts_467;
  wire [63:0] regOuts_468;
  wire [63:0] regOuts_469;
  wire [63:0] regOuts_470;
  wire [63:0] regOuts_471;
  wire [63:0] regOuts_472;
  wire [63:0] regOuts_473;
  wire [63:0] regOuts_474;
  wire [63:0] regOuts_475;
  wire [63:0] regOuts_476;
  wire [63:0] regOuts_477;
  wire [63:0] regOuts_478;
  wire [63:0] regOuts_479;
  wire [63:0] regOuts_480;
  wire [63:0] regOuts_481;
  wire [63:0] regOuts_482;
  wire [63:0] regOuts_483;
  wire [63:0] regOuts_484;
  wire [63:0] regOuts_485;
  wire [63:0] regOuts_486;
  wire [63:0] regOuts_487;
  wire [63:0] regOuts_488;
  wire [63:0] regOuts_489;
  wire [63:0] regOuts_490;
  wire [63:0] regOuts_491;
  wire [63:0] regOuts_492;
  wire [63:0] regOuts_493;
  wire [63:0] regOuts_494;
  wire [63:0] regOuts_495;
  wire [63:0] regOuts_496;
  wire [63:0] regOuts_497;
  wire [63:0] regOuts_498;
  wire [63:0] regOuts_499;
  wire [63:0] regOuts_500;
  wire [63:0] regOuts_501;
  wire [63:0] regOuts_502;
  wire [63:0] regOuts_503;
  wire [63:0] regOuts_504;
  wire [63:0] _T_5082_0;
  wire [63:0] _T_5082_1;
  wire [63:0] _T_5082_2;
  wire [63:0] _T_5082_3;
  FF_26 regs_0 (
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_init(regs_0_io_init),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FF_26 regs_1 (
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_init(regs_1_io_init),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FF_26 regs_2 (
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_init(regs_2_io_init),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FF_26 regs_3 (
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_init(regs_3_io_init),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FF_26 regs_4 (
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_init(regs_4_io_init),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FF_26 regs_5 (
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_init(regs_5_io_init),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FF_26 regs_6 (
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_init(regs_6_io_init),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FF_26 regs_7 (
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_init(regs_7_io_init),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FF_26 regs_8 (
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_init(regs_8_io_init),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FF_26 regs_9 (
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_init(regs_9_io_init),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FF_26 regs_10 (
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_init(regs_10_io_init),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FF_26 regs_11 (
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_init(regs_11_io_init),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FF_26 regs_12 (
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_init(regs_12_io_init),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FF_26 regs_13 (
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_init(regs_13_io_init),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FF_26 regs_14 (
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_init(regs_14_io_init),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FF_26 regs_15 (
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_init(regs_15_io_init),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FF_26 regs_16 (
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_init(regs_16_io_init),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FF_26 regs_17 (
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_init(regs_17_io_init),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FF_26 regs_18 (
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_init(regs_18_io_init),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FF_26 regs_19 (
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_init(regs_19_io_init),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FF_26 regs_20 (
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_init(regs_20_io_init),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FF_26 regs_21 (
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_init(regs_21_io_init),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FF_26 regs_22 (
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_init(regs_22_io_init),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FF_26 regs_23 (
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_init(regs_23_io_init),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FF_26 regs_24 (
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_init(regs_24_io_init),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FF_26 regs_25 (
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_init(regs_25_io_init),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FF_26 regs_26 (
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_init(regs_26_io_init),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FF_26 regs_27 (
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_init(regs_27_io_init),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FF_26 regs_28 (
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_init(regs_28_io_init),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FF_26 regs_29 (
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_init(regs_29_io_init),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FF_26 regs_30 (
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_init(regs_30_io_init),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FF_26 regs_31 (
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_init(regs_31_io_init),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FF_26 regs_32 (
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_init(regs_32_io_init),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FF_26 regs_33 (
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_init(regs_33_io_init),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FF_26 regs_34 (
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_init(regs_34_io_init),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FF_26 regs_35 (
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_init(regs_35_io_init),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FF_26 regs_36 (
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_init(regs_36_io_init),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FF_26 regs_37 (
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_init(regs_37_io_init),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FF_26 regs_38 (
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_init(regs_38_io_init),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FF_26 regs_39 (
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_init(regs_39_io_init),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FF_26 regs_40 (
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_init(regs_40_io_init),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FF_26 regs_41 (
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_init(regs_41_io_init),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FF_26 regs_42 (
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_init(regs_42_io_init),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FF_26 regs_43 (
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_init(regs_43_io_init),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FF_26 regs_44 (
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_init(regs_44_io_init),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FF_26 regs_45 (
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_init(regs_45_io_init),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FF_26 regs_46 (
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_init(regs_46_io_init),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FF_26 regs_47 (
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_init(regs_47_io_init),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FF_26 regs_48 (
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_init(regs_48_io_init),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FF_26 regs_49 (
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_init(regs_49_io_init),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FF_26 regs_50 (
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_init(regs_50_io_init),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FF_26 regs_51 (
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_init(regs_51_io_init),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FF_26 regs_52 (
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_init(regs_52_io_init),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FF_26 regs_53 (
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_init(regs_53_io_init),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FF_26 regs_54 (
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_init(regs_54_io_init),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FF_26 regs_55 (
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_init(regs_55_io_init),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FF_26 regs_56 (
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_init(regs_56_io_init),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FF_26 regs_57 (
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_init(regs_57_io_init),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FF_26 regs_58 (
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_init(regs_58_io_init),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FF_26 regs_59 (
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_init(regs_59_io_init),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FF_26 regs_60 (
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_init(regs_60_io_init),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FF_26 regs_61 (
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_init(regs_61_io_init),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FF_26 regs_62 (
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_init(regs_62_io_init),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FF_26 regs_63 (
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_init(regs_63_io_init),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FF_26 regs_64 (
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_init(regs_64_io_init),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FF_26 regs_65 (
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_init(regs_65_io_init),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FF_26 regs_66 (
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_init(regs_66_io_init),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FF_26 regs_67 (
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_init(regs_67_io_init),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FF_26 regs_68 (
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_init(regs_68_io_init),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FF_26 regs_69 (
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_init(regs_69_io_init),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FF_26 regs_70 (
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_init(regs_70_io_init),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FF_26 regs_71 (
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_init(regs_71_io_init),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FF_26 regs_72 (
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_init(regs_72_io_init),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FF_26 regs_73 (
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_init(regs_73_io_init),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FF_26 regs_74 (
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_init(regs_74_io_init),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FF_26 regs_75 (
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_init(regs_75_io_init),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FF_26 regs_76 (
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_init(regs_76_io_init),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FF_26 regs_77 (
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_init(regs_77_io_init),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FF_26 regs_78 (
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_init(regs_78_io_init),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FF_26 regs_79 (
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_init(regs_79_io_init),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FF_26 regs_80 (
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_init(regs_80_io_init),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FF_26 regs_81 (
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_init(regs_81_io_init),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FF_26 regs_82 (
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_init(regs_82_io_init),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FF_26 regs_83 (
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_init(regs_83_io_init),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FF_26 regs_84 (
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_init(regs_84_io_init),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FF_26 regs_85 (
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_init(regs_85_io_init),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FF_26 regs_86 (
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_init(regs_86_io_init),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FF_26 regs_87 (
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_init(regs_87_io_init),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FF_26 regs_88 (
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_init(regs_88_io_init),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FF_26 regs_89 (
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_init(regs_89_io_init),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FF_26 regs_90 (
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_init(regs_90_io_init),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FF_26 regs_91 (
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_init(regs_91_io_init),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FF_26 regs_92 (
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_init(regs_92_io_init),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FF_26 regs_93 (
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_init(regs_93_io_init),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FF_26 regs_94 (
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_init(regs_94_io_init),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FF_26 regs_95 (
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_init(regs_95_io_init),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FF_26 regs_96 (
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_init(regs_96_io_init),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FF_26 regs_97 (
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_init(regs_97_io_init),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FF_26 regs_98 (
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_init(regs_98_io_init),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FF_26 regs_99 (
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_init(regs_99_io_init),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FF_26 regs_100 (
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_init(regs_100_io_init),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FF_26 regs_101 (
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_init(regs_101_io_init),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FF_26 regs_102 (
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_init(regs_102_io_init),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FF_26 regs_103 (
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_init(regs_103_io_init),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FF_26 regs_104 (
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_init(regs_104_io_init),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FF_26 regs_105 (
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_init(regs_105_io_init),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FF_26 regs_106 (
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_init(regs_106_io_init),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FF_26 regs_107 (
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_init(regs_107_io_init),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FF_26 regs_108 (
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_init(regs_108_io_init),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FF_26 regs_109 (
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_init(regs_109_io_init),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FF_26 regs_110 (
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_init(regs_110_io_init),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FF_26 regs_111 (
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_init(regs_111_io_init),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FF_26 regs_112 (
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_init(regs_112_io_init),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FF_26 regs_113 (
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_init(regs_113_io_init),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FF_26 regs_114 (
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_init(regs_114_io_init),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FF_26 regs_115 (
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_init(regs_115_io_init),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FF_26 regs_116 (
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_init(regs_116_io_init),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FF_26 regs_117 (
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_init(regs_117_io_init),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FF_26 regs_118 (
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_init(regs_118_io_init),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FF_26 regs_119 (
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_init(regs_119_io_init),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FF_26 regs_120 (
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_init(regs_120_io_init),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FF_26 regs_121 (
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_init(regs_121_io_init),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FF_26 regs_122 (
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_init(regs_122_io_init),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FF_26 regs_123 (
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_init(regs_123_io_init),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FF_26 regs_124 (
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_init(regs_124_io_init),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FF_26 regs_125 (
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_init(regs_125_io_init),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FF_26 regs_126 (
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_init(regs_126_io_init),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FF_26 regs_127 (
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_init(regs_127_io_init),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FF_26 regs_128 (
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_init(regs_128_io_init),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FF_26 regs_129 (
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_init(regs_129_io_init),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FF_26 regs_130 (
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_init(regs_130_io_init),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FF_26 regs_131 (
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_init(regs_131_io_init),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FF_26 regs_132 (
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_init(regs_132_io_init),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FF_26 regs_133 (
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_init(regs_133_io_init),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FF_26 regs_134 (
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_init(regs_134_io_init),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FF_26 regs_135 (
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_init(regs_135_io_init),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FF_26 regs_136 (
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_init(regs_136_io_init),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FF_26 regs_137 (
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_init(regs_137_io_init),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FF_26 regs_138 (
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_init(regs_138_io_init),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FF_26 regs_139 (
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_init(regs_139_io_init),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FF_26 regs_140 (
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_init(regs_140_io_init),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FF_26 regs_141 (
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_init(regs_141_io_init),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FF_26 regs_142 (
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_init(regs_142_io_init),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FF_26 regs_143 (
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_init(regs_143_io_init),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FF_26 regs_144 (
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_init(regs_144_io_init),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FF_26 regs_145 (
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_init(regs_145_io_init),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FF_26 regs_146 (
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_init(regs_146_io_init),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FF_26 regs_147 (
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_init(regs_147_io_init),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FF_26 regs_148 (
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_init(regs_148_io_init),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FF_26 regs_149 (
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_init(regs_149_io_init),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FF_26 regs_150 (
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_init(regs_150_io_init),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FF_26 regs_151 (
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_init(regs_151_io_init),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FF_26 regs_152 (
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_init(regs_152_io_init),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FF_26 regs_153 (
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_init(regs_153_io_init),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FF_26 regs_154 (
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_init(regs_154_io_init),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FF_26 regs_155 (
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_init(regs_155_io_init),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FF_26 regs_156 (
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_init(regs_156_io_init),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FF_26 regs_157 (
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_init(regs_157_io_init),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FF_26 regs_158 (
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_init(regs_158_io_init),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FF_26 regs_159 (
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_init(regs_159_io_init),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FF_26 regs_160 (
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_init(regs_160_io_init),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FF_26 regs_161 (
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_init(regs_161_io_init),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FF_26 regs_162 (
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_init(regs_162_io_init),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FF_26 regs_163 (
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_init(regs_163_io_init),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FF_26 regs_164 (
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_init(regs_164_io_init),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FF_26 regs_165 (
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_init(regs_165_io_init),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FF_26 regs_166 (
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_init(regs_166_io_init),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FF_26 regs_167 (
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_init(regs_167_io_init),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FF_26 regs_168 (
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_init(regs_168_io_init),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FF_26 regs_169 (
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_init(regs_169_io_init),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FF_26 regs_170 (
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_init(regs_170_io_init),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FF_26 regs_171 (
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_init(regs_171_io_init),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FF_26 regs_172 (
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_init(regs_172_io_init),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FF_26 regs_173 (
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_init(regs_173_io_init),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FF_26 regs_174 (
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_init(regs_174_io_init),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FF_26 regs_175 (
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_init(regs_175_io_init),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FF_26 regs_176 (
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_init(regs_176_io_init),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FF_26 regs_177 (
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_init(regs_177_io_init),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FF_26 regs_178 (
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_init(regs_178_io_init),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FF_26 regs_179 (
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_init(regs_179_io_init),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FF_26 regs_180 (
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_init(regs_180_io_init),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FF_26 regs_181 (
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_init(regs_181_io_init),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FF_26 regs_182 (
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_init(regs_182_io_init),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FF_26 regs_183 (
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_init(regs_183_io_init),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FF_26 regs_184 (
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_init(regs_184_io_init),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FF_26 regs_185 (
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_init(regs_185_io_init),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FF_26 regs_186 (
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_init(regs_186_io_init),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FF_26 regs_187 (
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_init(regs_187_io_init),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FF_26 regs_188 (
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_init(regs_188_io_init),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FF_26 regs_189 (
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_init(regs_189_io_init),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FF_26 regs_190 (
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_init(regs_190_io_init),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FF_26 regs_191 (
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_init(regs_191_io_init),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FF_26 regs_192 (
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_init(regs_192_io_init),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FF_26 regs_193 (
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_init(regs_193_io_init),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FF_26 regs_194 (
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_init(regs_194_io_init),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FF_26 regs_195 (
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_init(regs_195_io_init),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FF_26 regs_196 (
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_init(regs_196_io_init),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FF_26 regs_197 (
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_init(regs_197_io_init),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FF_26 regs_198 (
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_init(regs_198_io_init),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FF_26 regs_199 (
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_init(regs_199_io_init),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FF_26 regs_200 (
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_init(regs_200_io_init),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FF_26 regs_201 (
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_init(regs_201_io_init),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FF_26 regs_202 (
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_init(regs_202_io_init),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FF_26 regs_203 (
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_init(regs_203_io_init),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FF_26 regs_204 (
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_init(regs_204_io_init),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FF_26 regs_205 (
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_init(regs_205_io_init),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FF_26 regs_206 (
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_init(regs_206_io_init),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FF_26 regs_207 (
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_init(regs_207_io_init),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FF_26 regs_208 (
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_init(regs_208_io_init),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FF_26 regs_209 (
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_init(regs_209_io_init),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FF_26 regs_210 (
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_init(regs_210_io_init),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FF_26 regs_211 (
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_init(regs_211_io_init),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FF_26 regs_212 (
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_init(regs_212_io_init),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FF_26 regs_213 (
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_init(regs_213_io_init),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FF_26 regs_214 (
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_init(regs_214_io_init),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FF_26 regs_215 (
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_init(regs_215_io_init),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FF_26 regs_216 (
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_init(regs_216_io_init),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FF_26 regs_217 (
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_init(regs_217_io_init),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FF_26 regs_218 (
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_init(regs_218_io_init),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FF_26 regs_219 (
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_init(regs_219_io_init),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FF_26 regs_220 (
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_init(regs_220_io_init),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FF_26 regs_221 (
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_init(regs_221_io_init),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FF_26 regs_222 (
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_init(regs_222_io_init),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FF_26 regs_223 (
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_init(regs_223_io_init),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FF_26 regs_224 (
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_init(regs_224_io_init),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FF_26 regs_225 (
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_init(regs_225_io_init),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FF_26 regs_226 (
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_init(regs_226_io_init),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FF_26 regs_227 (
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_init(regs_227_io_init),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FF_26 regs_228 (
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_init(regs_228_io_init),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FF_26 regs_229 (
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_init(regs_229_io_init),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FF_26 regs_230 (
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_init(regs_230_io_init),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FF_26 regs_231 (
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_init(regs_231_io_init),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FF_26 regs_232 (
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_init(regs_232_io_init),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FF_26 regs_233 (
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_init(regs_233_io_init),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FF_26 regs_234 (
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_init(regs_234_io_init),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FF_26 regs_235 (
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_init(regs_235_io_init),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FF_26 regs_236 (
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_init(regs_236_io_init),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FF_26 regs_237 (
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_init(regs_237_io_init),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FF_26 regs_238 (
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_init(regs_238_io_init),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FF_26 regs_239 (
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_init(regs_239_io_init),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FF_26 regs_240 (
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_init(regs_240_io_init),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FF_26 regs_241 (
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_init(regs_241_io_init),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FF_26 regs_242 (
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_init(regs_242_io_init),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FF_26 regs_243 (
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_init(regs_243_io_init),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FF_26 regs_244 (
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_init(regs_244_io_init),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FF_26 regs_245 (
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_init(regs_245_io_init),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FF_26 regs_246 (
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_init(regs_246_io_init),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FF_26 regs_247 (
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_init(regs_247_io_init),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FF_26 regs_248 (
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_init(regs_248_io_init),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FF_26 regs_249 (
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_init(regs_249_io_init),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FF_26 regs_250 (
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_init(regs_250_io_init),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FF_26 regs_251 (
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_init(regs_251_io_init),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FF_26 regs_252 (
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_init(regs_252_io_init),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FF_26 regs_253 (
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_init(regs_253_io_init),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FF_26 regs_254 (
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_init(regs_254_io_init),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FF_26 regs_255 (
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_init(regs_255_io_init),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FF_26 regs_256 (
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_init(regs_256_io_init),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FF_26 regs_257 (
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_init(regs_257_io_init),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FF_26 regs_258 (
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_init(regs_258_io_init),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FF_26 regs_259 (
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_init(regs_259_io_init),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FF_26 regs_260 (
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_init(regs_260_io_init),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FF_26 regs_261 (
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_init(regs_261_io_init),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FF_26 regs_262 (
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_init(regs_262_io_init),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FF_26 regs_263 (
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_init(regs_263_io_init),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FF_26 regs_264 (
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_init(regs_264_io_init),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FF_26 regs_265 (
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_init(regs_265_io_init),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FF_26 regs_266 (
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_init(regs_266_io_init),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FF_26 regs_267 (
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_init(regs_267_io_init),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FF_26 regs_268 (
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_init(regs_268_io_init),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FF_26 regs_269 (
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_init(regs_269_io_init),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FF_26 regs_270 (
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_init(regs_270_io_init),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FF_26 regs_271 (
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_init(regs_271_io_init),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FF_26 regs_272 (
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_init(regs_272_io_init),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FF_26 regs_273 (
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_init(regs_273_io_init),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FF_26 regs_274 (
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_init(regs_274_io_init),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FF_26 regs_275 (
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_init(regs_275_io_init),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FF_26 regs_276 (
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_init(regs_276_io_init),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FF_26 regs_277 (
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_init(regs_277_io_init),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FF_26 regs_278 (
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_init(regs_278_io_init),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FF_26 regs_279 (
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_init(regs_279_io_init),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FF_26 regs_280 (
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_init(regs_280_io_init),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FF_26 regs_281 (
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_init(regs_281_io_init),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FF_26 regs_282 (
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_init(regs_282_io_init),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FF_26 regs_283 (
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_init(regs_283_io_init),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FF_26 regs_284 (
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_init(regs_284_io_init),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FF_26 regs_285 (
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_init(regs_285_io_init),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FF_26 regs_286 (
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_init(regs_286_io_init),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FF_26 regs_287 (
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_init(regs_287_io_init),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FF_26 regs_288 (
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_init(regs_288_io_init),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FF_26 regs_289 (
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_init(regs_289_io_init),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FF_26 regs_290 (
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_init(regs_290_io_init),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FF_26 regs_291 (
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_init(regs_291_io_init),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FF_26 regs_292 (
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_init(regs_292_io_init),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FF_26 regs_293 (
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_init(regs_293_io_init),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FF_26 regs_294 (
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_init(regs_294_io_init),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FF_26 regs_295 (
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_init(regs_295_io_init),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FF_26 regs_296 (
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_init(regs_296_io_init),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FF_26 regs_297 (
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_init(regs_297_io_init),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FF_26 regs_298 (
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_init(regs_298_io_init),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FF_26 regs_299 (
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_init(regs_299_io_init),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FF_26 regs_300 (
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_init(regs_300_io_init),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FF_26 regs_301 (
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_init(regs_301_io_init),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FF_26 regs_302 (
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_init(regs_302_io_init),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FF_26 regs_303 (
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_init(regs_303_io_init),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FF_26 regs_304 (
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_init(regs_304_io_init),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FF_26 regs_305 (
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_init(regs_305_io_init),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FF_26 regs_306 (
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_init(regs_306_io_init),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FF_26 regs_307 (
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_init(regs_307_io_init),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FF_26 regs_308 (
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_init(regs_308_io_init),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FF_26 regs_309 (
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_init(regs_309_io_init),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FF_26 regs_310 (
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_init(regs_310_io_init),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FF_26 regs_311 (
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_init(regs_311_io_init),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FF_26 regs_312 (
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_init(regs_312_io_init),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FF_26 regs_313 (
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_init(regs_313_io_init),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FF_26 regs_314 (
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_init(regs_314_io_init),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FF_26 regs_315 (
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_init(regs_315_io_init),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FF_26 regs_316 (
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_init(regs_316_io_init),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FF_26 regs_317 (
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_init(regs_317_io_init),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FF_26 regs_318 (
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_init(regs_318_io_init),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FF_26 regs_319 (
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_init(regs_319_io_init),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FF_26 regs_320 (
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_init(regs_320_io_init),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FF_26 regs_321 (
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_init(regs_321_io_init),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FF_26 regs_322 (
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_init(regs_322_io_init),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FF_26 regs_323 (
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_init(regs_323_io_init),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FF_26 regs_324 (
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_init(regs_324_io_init),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FF_26 regs_325 (
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_init(regs_325_io_init),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FF_26 regs_326 (
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_init(regs_326_io_init),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FF_26 regs_327 (
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_init(regs_327_io_init),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FF_26 regs_328 (
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_init(regs_328_io_init),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FF_26 regs_329 (
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_init(regs_329_io_init),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FF_26 regs_330 (
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_init(regs_330_io_init),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FF_26 regs_331 (
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_init(regs_331_io_init),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FF_26 regs_332 (
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_init(regs_332_io_init),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FF_26 regs_333 (
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_init(regs_333_io_init),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FF_26 regs_334 (
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_init(regs_334_io_init),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FF_26 regs_335 (
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_init(regs_335_io_init),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FF_26 regs_336 (
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_init(regs_336_io_init),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FF_26 regs_337 (
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_init(regs_337_io_init),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FF_26 regs_338 (
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_init(regs_338_io_init),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FF_26 regs_339 (
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_init(regs_339_io_init),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FF_26 regs_340 (
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_init(regs_340_io_init),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FF_26 regs_341 (
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_init(regs_341_io_init),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FF_26 regs_342 (
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_init(regs_342_io_init),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FF_26 regs_343 (
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_init(regs_343_io_init),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FF_26 regs_344 (
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_init(regs_344_io_init),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FF_26 regs_345 (
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_init(regs_345_io_init),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FF_26 regs_346 (
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_init(regs_346_io_init),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FF_26 regs_347 (
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_init(regs_347_io_init),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FF_26 regs_348 (
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_init(regs_348_io_init),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FF_26 regs_349 (
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_init(regs_349_io_init),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FF_26 regs_350 (
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_init(regs_350_io_init),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FF_26 regs_351 (
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_init(regs_351_io_init),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FF_26 regs_352 (
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_init(regs_352_io_init),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FF_26 regs_353 (
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_init(regs_353_io_init),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FF_26 regs_354 (
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_init(regs_354_io_init),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FF_26 regs_355 (
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_init(regs_355_io_init),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FF_26 regs_356 (
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_init(regs_356_io_init),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FF_26 regs_357 (
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_init(regs_357_io_init),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FF_26 regs_358 (
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_init(regs_358_io_init),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FF_26 regs_359 (
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_init(regs_359_io_init),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FF_26 regs_360 (
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_init(regs_360_io_init),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FF_26 regs_361 (
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_init(regs_361_io_init),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FF_26 regs_362 (
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_init(regs_362_io_init),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FF_26 regs_363 (
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_init(regs_363_io_init),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FF_26 regs_364 (
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_init(regs_364_io_init),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FF_26 regs_365 (
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_init(regs_365_io_init),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FF_26 regs_366 (
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_init(regs_366_io_init),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FF_26 regs_367 (
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_init(regs_367_io_init),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FF_26 regs_368 (
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_init(regs_368_io_init),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FF_26 regs_369 (
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_init(regs_369_io_init),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FF_26 regs_370 (
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_init(regs_370_io_init),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FF_26 regs_371 (
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_init(regs_371_io_init),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FF_26 regs_372 (
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_init(regs_372_io_init),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FF_26 regs_373 (
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_init(regs_373_io_init),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FF_26 regs_374 (
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_init(regs_374_io_init),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FF_26 regs_375 (
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_init(regs_375_io_init),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FF_26 regs_376 (
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_init(regs_376_io_init),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FF_26 regs_377 (
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_init(regs_377_io_init),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FF_26 regs_378 (
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_init(regs_378_io_init),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FF_26 regs_379 (
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_init(regs_379_io_init),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FF_26 regs_380 (
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_init(regs_380_io_init),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FF_26 regs_381 (
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_init(regs_381_io_init),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FF_26 regs_382 (
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_init(regs_382_io_init),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FF_26 regs_383 (
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_init(regs_383_io_init),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FF_26 regs_384 (
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_init(regs_384_io_init),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FF_26 regs_385 (
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_init(regs_385_io_init),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FF_26 regs_386 (
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_init(regs_386_io_init),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FF_26 regs_387 (
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_init(regs_387_io_init),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FF_26 regs_388 (
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_init(regs_388_io_init),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FF_26 regs_389 (
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_init(regs_389_io_init),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FF_26 regs_390 (
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_init(regs_390_io_init),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FF_26 regs_391 (
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_init(regs_391_io_init),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FF_26 regs_392 (
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_init(regs_392_io_init),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FF_26 regs_393 (
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_init(regs_393_io_init),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FF_26 regs_394 (
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_init(regs_394_io_init),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FF_26 regs_395 (
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_init(regs_395_io_init),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FF_26 regs_396 (
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_init(regs_396_io_init),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FF_26 regs_397 (
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_init(regs_397_io_init),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FF_26 regs_398 (
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_init(regs_398_io_init),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FF_26 regs_399 (
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_init(regs_399_io_init),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FF_26 regs_400 (
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_init(regs_400_io_init),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FF_26 regs_401 (
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_init(regs_401_io_init),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FF_26 regs_402 (
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_init(regs_402_io_init),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FF_26 regs_403 (
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_init(regs_403_io_init),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FF_26 regs_404 (
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_init(regs_404_io_init),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FF_26 regs_405 (
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_init(regs_405_io_init),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FF_26 regs_406 (
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_init(regs_406_io_init),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FF_26 regs_407 (
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_init(regs_407_io_init),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FF_26 regs_408 (
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_init(regs_408_io_init),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FF_26 regs_409 (
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_init(regs_409_io_init),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FF_26 regs_410 (
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_init(regs_410_io_init),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FF_26 regs_411 (
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_init(regs_411_io_init),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FF_26 regs_412 (
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_init(regs_412_io_init),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FF_26 regs_413 (
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_init(regs_413_io_init),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FF_26 regs_414 (
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_init(regs_414_io_init),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FF_26 regs_415 (
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_init(regs_415_io_init),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FF_26 regs_416 (
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_init(regs_416_io_init),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FF_26 regs_417 (
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_init(regs_417_io_init),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FF_26 regs_418 (
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_init(regs_418_io_init),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FF_26 regs_419 (
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_init(regs_419_io_init),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FF_26 regs_420 (
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_init(regs_420_io_init),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FF_26 regs_421 (
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_init(regs_421_io_init),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FF_26 regs_422 (
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_init(regs_422_io_init),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FF_26 regs_423 (
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_init(regs_423_io_init),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FF_26 regs_424 (
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_init(regs_424_io_init),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FF_26 regs_425 (
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_init(regs_425_io_init),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FF_26 regs_426 (
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_init(regs_426_io_init),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FF_26 regs_427 (
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_init(regs_427_io_init),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FF_26 regs_428 (
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_init(regs_428_io_init),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FF_26 regs_429 (
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_init(regs_429_io_init),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FF_26 regs_430 (
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_init(regs_430_io_init),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FF_26 regs_431 (
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_init(regs_431_io_init),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FF_26 regs_432 (
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_init(regs_432_io_init),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FF_26 regs_433 (
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_init(regs_433_io_init),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FF_26 regs_434 (
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_init(regs_434_io_init),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FF_26 regs_435 (
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_init(regs_435_io_init),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FF_26 regs_436 (
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_init(regs_436_io_init),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FF_26 regs_437 (
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_init(regs_437_io_init),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FF_26 regs_438 (
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_init(regs_438_io_init),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FF_26 regs_439 (
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_init(regs_439_io_init),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FF_26 regs_440 (
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_init(regs_440_io_init),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FF_26 regs_441 (
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_init(regs_441_io_init),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FF_26 regs_442 (
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_init(regs_442_io_init),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FF_26 regs_443 (
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_init(regs_443_io_init),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FF_26 regs_444 (
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_init(regs_444_io_init),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FF_26 regs_445 (
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_init(regs_445_io_init),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FF_26 regs_446 (
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_init(regs_446_io_init),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FF_26 regs_447 (
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_init(regs_447_io_init),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FF_26 regs_448 (
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_init(regs_448_io_init),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FF_26 regs_449 (
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_init(regs_449_io_init),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FF_26 regs_450 (
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_init(regs_450_io_init),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FF_26 regs_451 (
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_init(regs_451_io_init),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FF_26 regs_452 (
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_init(regs_452_io_init),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FF_26 regs_453 (
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_init(regs_453_io_init),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FF_26 regs_454 (
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_init(regs_454_io_init),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FF_26 regs_455 (
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_init(regs_455_io_init),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FF_26 regs_456 (
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_init(regs_456_io_init),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FF_26 regs_457 (
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_init(regs_457_io_init),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FF_26 regs_458 (
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_init(regs_458_io_init),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FF_26 regs_459 (
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_init(regs_459_io_init),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FF_26 regs_460 (
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_init(regs_460_io_init),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FF_26 regs_461 (
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_init(regs_461_io_init),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FF_26 regs_462 (
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_init(regs_462_io_init),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FF_26 regs_463 (
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_init(regs_463_io_init),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FF_26 regs_464 (
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_init(regs_464_io_init),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FF_26 regs_465 (
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_init(regs_465_io_init),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FF_26 regs_466 (
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_init(regs_466_io_init),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FF_26 regs_467 (
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_init(regs_467_io_init),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FF_26 regs_468 (
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_init(regs_468_io_init),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FF_26 regs_469 (
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_init(regs_469_io_init),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FF_26 regs_470 (
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_init(regs_470_io_init),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FF_26 regs_471 (
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_init(regs_471_io_init),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FF_26 regs_472 (
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_init(regs_472_io_init),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FF_26 regs_473 (
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_init(regs_473_io_init),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FF_26 regs_474 (
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_init(regs_474_io_init),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FF_26 regs_475 (
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_init(regs_475_io_init),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FF_26 regs_476 (
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_init(regs_476_io_init),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FF_26 regs_477 (
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_init(regs_477_io_init),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FF_26 regs_478 (
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_init(regs_478_io_init),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FF_26 regs_479 (
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_init(regs_479_io_init),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FF_26 regs_480 (
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_init(regs_480_io_init),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FF_26 regs_481 (
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_init(regs_481_io_init),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FF_26 regs_482 (
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_init(regs_482_io_init),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FF_26 regs_483 (
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_init(regs_483_io_init),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FF_26 regs_484 (
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_init(regs_484_io_init),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FF_26 regs_485 (
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_init(regs_485_io_init),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FF_26 regs_486 (
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_init(regs_486_io_init),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FF_26 regs_487 (
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_init(regs_487_io_init),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FF_26 regs_488 (
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_init(regs_488_io_init),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FF_26 regs_489 (
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_init(regs_489_io_init),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FF_26 regs_490 (
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_init(regs_490_io_init),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FF_26 regs_491 (
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_init(regs_491_io_init),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FF_26 regs_492 (
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_init(regs_492_io_init),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FF_26 regs_493 (
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_init(regs_493_io_init),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FF_26 regs_494 (
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_init(regs_494_io_init),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FF_26 regs_495 (
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_init(regs_495_io_init),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FF_26 regs_496 (
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_init(regs_496_io_init),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FF_26 regs_497 (
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_init(regs_497_io_init),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FF_26 regs_498 (
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_init(regs_498_io_init),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FF_26 regs_499 (
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_init(regs_499_io_init),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FF_26 regs_500 (
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_init(regs_500_io_init),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FF_26 regs_501 (
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_init(regs_501_io_init),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FF_26 regs_502 (
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_init(regs_502_io_init),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  FF_26 regs_503 (
    .clock(regs_503_clock),
    .reset(regs_503_reset),
    .io_in(regs_503_io_in),
    .io_init(regs_503_io_init),
    .io_out(regs_503_io_out),
    .io_enable(regs_503_io_enable)
  );
  FF_26 regs_504 (
    .clock(regs_504_clock),
    .reset(regs_504_reset),
    .io_in(regs_504_io_in),
    .io_init(regs_504_io_init),
    .io_out(regs_504_io_out),
    .io_enable(regs_504_io_enable)
  );
  MuxN_16 rport (
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_ins_503(rport_io_ins_503),
    .io_ins_504(rport_io_ins_504),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_1542 = io_waddr == 9'h0;
  assign _T_1543 = io_wen & _T_1542;
  assign _T_1546 = io_waddr == 9'h1;
  assign _T_1547 = io_wen & _T_1546;
  assign _T_1551 = _T_1547 ? _T_1547 : io_argOuts_0_valid;
  assign _T_1555 = _T_1547 ? io_wdata : io_argOuts_0_bits;
  assign _T_1558 = io_waddr == 9'h2;
  assign _T_1559 = io_wen & _T_1558;
  assign _T_1562 = io_waddr == 9'h3;
  assign _T_1563 = io_wen & _T_1562;
  assign _T_1566 = io_waddr == 9'h4;
  assign _T_1567 = io_wen & _T_1566;
  assign _T_1568 = io_argOuts_1_valid | _T_1567;
  assign _T_1569 = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata;
  assign io_rdata = rport_io_out;
  assign io_argIns_0 = _T_5082_0;
  assign io_argIns_1 = _T_5082_1;
  assign io_argIns_2 = _T_5082_2;
  assign io_argIns_3 = _T_5082_3;
  assign regs_0_io_in = io_wdata;
  assign regs_0_io_init = 64'h0;
  assign regs_0_io_enable = _T_1543;
  assign regs_0_clock = clock;
  assign regs_0_reset = reset;
  assign regs_1_io_in = _T_1555;
  assign regs_1_io_init = 64'h0;
  assign regs_1_io_enable = _T_1551;
  assign regs_1_clock = clock;
  assign regs_1_reset = reset;
  assign regs_2_io_in = io_wdata;
  assign regs_2_io_init = 64'h0;
  assign regs_2_io_enable = _T_1559;
  assign regs_2_clock = clock;
  assign regs_2_reset = reset;
  assign regs_3_io_in = io_wdata;
  assign regs_3_io_init = 64'h0;
  assign regs_3_io_enable = _T_1563;
  assign regs_3_clock = clock;
  assign regs_3_reset = reset;
  assign regs_4_io_in = _T_1569;
  assign regs_4_io_init = 64'h0;
  assign regs_4_io_enable = _T_1568;
  assign regs_4_clock = clock;
  assign regs_4_reset = reset;
  assign regs_5_io_in = io_argOuts_2_bits;
  assign regs_5_io_init = 64'h0;
  assign regs_5_io_enable = 1'h1;
  assign regs_5_clock = clock;
  assign regs_5_reset = reset;
  assign regs_6_io_in = io_argOuts_3_bits;
  assign regs_6_io_init = 64'h0;
  assign regs_6_io_enable = 1'h1;
  assign regs_6_clock = clock;
  assign regs_6_reset = reset;
  assign regs_7_io_in = io_argOuts_4_bits;
  assign regs_7_io_init = 64'h0;
  assign regs_7_io_enable = 1'h1;
  assign regs_7_clock = clock;
  assign regs_7_reset = reset;
  assign regs_8_io_in = io_argOuts_5_bits;
  assign regs_8_io_init = 64'h0;
  assign regs_8_io_enable = 1'h1;
  assign regs_8_clock = clock;
  assign regs_8_reset = reset;
  assign regs_9_io_in = io_argOuts_6_bits;
  assign regs_9_io_init = 64'h0;
  assign regs_9_io_enable = 1'h1;
  assign regs_9_clock = clock;
  assign regs_9_reset = reset;
  assign regs_10_io_in = io_argOuts_7_bits;
  assign regs_10_io_init = 64'h0;
  assign regs_10_io_enable = 1'h1;
  assign regs_10_clock = clock;
  assign regs_10_reset = reset;
  assign regs_11_io_in = io_argOuts_8_bits;
  assign regs_11_io_init = 64'h0;
  assign regs_11_io_enable = 1'h1;
  assign regs_11_clock = clock;
  assign regs_11_reset = reset;
  assign regs_12_io_in = io_argOuts_9_bits;
  assign regs_12_io_init = 64'h0;
  assign regs_12_io_enable = 1'h1;
  assign regs_12_clock = clock;
  assign regs_12_reset = reset;
  assign regs_13_io_in = io_argOuts_10_bits;
  assign regs_13_io_init = 64'h0;
  assign regs_13_io_enable = 1'h1;
  assign regs_13_clock = clock;
  assign regs_13_reset = reset;
  assign regs_14_io_in = io_argOuts_11_bits;
  assign regs_14_io_init = 64'h0;
  assign regs_14_io_enable = 1'h1;
  assign regs_14_clock = clock;
  assign regs_14_reset = reset;
  assign regs_15_io_in = io_argOuts_12_bits;
  assign regs_15_io_init = 64'h0;
  assign regs_15_io_enable = 1'h1;
  assign regs_15_clock = clock;
  assign regs_15_reset = reset;
  assign regs_16_io_in = io_argOuts_13_bits;
  assign regs_16_io_init = 64'h0;
  assign regs_16_io_enable = 1'h1;
  assign regs_16_clock = clock;
  assign regs_16_reset = reset;
  assign regs_17_io_in = io_argOuts_14_bits;
  assign regs_17_io_init = 64'h0;
  assign regs_17_io_enable = 1'h1;
  assign regs_17_clock = clock;
  assign regs_17_reset = reset;
  assign regs_18_io_in = io_argOuts_15_bits;
  assign regs_18_io_init = 64'h0;
  assign regs_18_io_enable = 1'h1;
  assign regs_18_clock = clock;
  assign regs_18_reset = reset;
  assign regs_19_io_in = io_argOuts_16_bits;
  assign regs_19_io_init = 64'h0;
  assign regs_19_io_enable = 1'h1;
  assign regs_19_clock = clock;
  assign regs_19_reset = reset;
  assign regs_20_io_in = io_argOuts_17_bits;
  assign regs_20_io_init = 64'h0;
  assign regs_20_io_enable = 1'h1;
  assign regs_20_clock = clock;
  assign regs_20_reset = reset;
  assign regs_21_io_in = io_argOuts_18_bits;
  assign regs_21_io_init = 64'h0;
  assign regs_21_io_enable = 1'h1;
  assign regs_21_clock = clock;
  assign regs_21_reset = reset;
  assign regs_22_io_in = io_argOuts_19_bits;
  assign regs_22_io_init = 64'h0;
  assign regs_22_io_enable = 1'h1;
  assign regs_22_clock = clock;
  assign regs_22_reset = reset;
  assign regs_23_io_in = io_argOuts_20_bits;
  assign regs_23_io_init = 64'h0;
  assign regs_23_io_enable = 1'h1;
  assign regs_23_clock = clock;
  assign regs_23_reset = reset;
  assign regs_24_io_in = io_argOuts_21_bits;
  assign regs_24_io_init = 64'h0;
  assign regs_24_io_enable = 1'h1;
  assign regs_24_clock = clock;
  assign regs_24_reset = reset;
  assign regs_25_io_in = io_argOuts_22_bits;
  assign regs_25_io_init = 64'h0;
  assign regs_25_io_enable = 1'h1;
  assign regs_25_clock = clock;
  assign regs_25_reset = reset;
  assign regs_26_io_in = io_argOuts_23_bits;
  assign regs_26_io_init = 64'h0;
  assign regs_26_io_enable = 1'h1;
  assign regs_26_clock = clock;
  assign regs_26_reset = reset;
  assign regs_27_io_in = io_argOuts_24_bits;
  assign regs_27_io_init = 64'h0;
  assign regs_27_io_enable = 1'h1;
  assign regs_27_clock = clock;
  assign regs_27_reset = reset;
  assign regs_28_io_in = io_argOuts_25_bits;
  assign regs_28_io_init = 64'h0;
  assign regs_28_io_enable = 1'h1;
  assign regs_28_clock = clock;
  assign regs_28_reset = reset;
  assign regs_29_io_in = io_argOuts_26_bits;
  assign regs_29_io_init = 64'h0;
  assign regs_29_io_enable = 1'h1;
  assign regs_29_clock = clock;
  assign regs_29_reset = reset;
  assign regs_30_io_in = io_argOuts_27_bits;
  assign regs_30_io_init = 64'h0;
  assign regs_30_io_enable = 1'h1;
  assign regs_30_clock = clock;
  assign regs_30_reset = reset;
  assign regs_31_io_in = io_argOuts_28_bits;
  assign regs_31_io_init = 64'h0;
  assign regs_31_io_enable = 1'h1;
  assign regs_31_clock = clock;
  assign regs_31_reset = reset;
  assign regs_32_io_in = io_argOuts_29_bits;
  assign regs_32_io_init = 64'h0;
  assign regs_32_io_enable = 1'h1;
  assign regs_32_clock = clock;
  assign regs_32_reset = reset;
  assign regs_33_io_in = io_argOuts_30_bits;
  assign regs_33_io_init = 64'h0;
  assign regs_33_io_enable = 1'h1;
  assign regs_33_clock = clock;
  assign regs_33_reset = reset;
  assign regs_34_io_in = io_argOuts_31_bits;
  assign regs_34_io_init = 64'h0;
  assign regs_34_io_enable = 1'h1;
  assign regs_34_clock = clock;
  assign regs_34_reset = reset;
  assign regs_35_io_in = io_argOuts_32_bits;
  assign regs_35_io_init = 64'h0;
  assign regs_35_io_enable = 1'h1;
  assign regs_35_clock = clock;
  assign regs_35_reset = reset;
  assign regs_36_io_in = io_argOuts_33_bits;
  assign regs_36_io_init = 64'h0;
  assign regs_36_io_enable = 1'h1;
  assign regs_36_clock = clock;
  assign regs_36_reset = reset;
  assign regs_37_io_in = io_argOuts_34_bits;
  assign regs_37_io_init = 64'h0;
  assign regs_37_io_enable = 1'h1;
  assign regs_37_clock = clock;
  assign regs_37_reset = reset;
  assign regs_38_io_in = io_argOuts_35_bits;
  assign regs_38_io_init = 64'h0;
  assign regs_38_io_enable = 1'h1;
  assign regs_38_clock = clock;
  assign regs_38_reset = reset;
  assign regs_39_io_in = io_argOuts_36_bits;
  assign regs_39_io_init = 64'h0;
  assign regs_39_io_enable = 1'h1;
  assign regs_39_clock = clock;
  assign regs_39_reset = reset;
  assign regs_40_io_in = io_argOuts_37_bits;
  assign regs_40_io_init = 64'h0;
  assign regs_40_io_enable = 1'h1;
  assign regs_40_clock = clock;
  assign regs_40_reset = reset;
  assign regs_41_io_in = io_argOuts_38_bits;
  assign regs_41_io_init = 64'h0;
  assign regs_41_io_enable = 1'h1;
  assign regs_41_clock = clock;
  assign regs_41_reset = reset;
  assign regs_42_io_in = io_argOuts_39_bits;
  assign regs_42_io_init = 64'h0;
  assign regs_42_io_enable = 1'h1;
  assign regs_42_clock = clock;
  assign regs_42_reset = reset;
  assign regs_43_io_in = io_argOuts_40_bits;
  assign regs_43_io_init = 64'h0;
  assign regs_43_io_enable = 1'h1;
  assign regs_43_clock = clock;
  assign regs_43_reset = reset;
  assign regs_44_io_in = io_argOuts_41_bits;
  assign regs_44_io_init = 64'h0;
  assign regs_44_io_enable = 1'h1;
  assign regs_44_clock = clock;
  assign regs_44_reset = reset;
  assign regs_45_io_in = io_argOuts_42_bits;
  assign regs_45_io_init = 64'h0;
  assign regs_45_io_enable = 1'h1;
  assign regs_45_clock = clock;
  assign regs_45_reset = reset;
  assign regs_46_io_in = io_argOuts_43_bits;
  assign regs_46_io_init = 64'h0;
  assign regs_46_io_enable = 1'h1;
  assign regs_46_clock = clock;
  assign regs_46_reset = reset;
  assign regs_47_io_in = io_argOuts_44_bits;
  assign regs_47_io_init = 64'h0;
  assign regs_47_io_enable = 1'h1;
  assign regs_47_clock = clock;
  assign regs_47_reset = reset;
  assign regs_48_io_in = io_argOuts_45_bits;
  assign regs_48_io_init = 64'h0;
  assign regs_48_io_enable = 1'h1;
  assign regs_48_clock = clock;
  assign regs_48_reset = reset;
  assign regs_49_io_in = io_argOuts_46_bits;
  assign regs_49_io_init = 64'h0;
  assign regs_49_io_enable = 1'h1;
  assign regs_49_clock = clock;
  assign regs_49_reset = reset;
  assign regs_50_io_in = io_argOuts_47_bits;
  assign regs_50_io_init = 64'h0;
  assign regs_50_io_enable = 1'h1;
  assign regs_50_clock = clock;
  assign regs_50_reset = reset;
  assign regs_51_io_in = io_argOuts_48_bits;
  assign regs_51_io_init = 64'h0;
  assign regs_51_io_enable = 1'h1;
  assign regs_51_clock = clock;
  assign regs_51_reset = reset;
  assign regs_52_io_in = io_argOuts_49_bits;
  assign regs_52_io_init = 64'h0;
  assign regs_52_io_enable = 1'h1;
  assign regs_52_clock = clock;
  assign regs_52_reset = reset;
  assign regs_53_io_in = io_argOuts_50_bits;
  assign regs_53_io_init = 64'h0;
  assign regs_53_io_enable = 1'h1;
  assign regs_53_clock = clock;
  assign regs_53_reset = reset;
  assign regs_54_io_in = io_argOuts_51_bits;
  assign regs_54_io_init = 64'h0;
  assign regs_54_io_enable = 1'h1;
  assign regs_54_clock = clock;
  assign regs_54_reset = reset;
  assign regs_55_io_in = io_argOuts_52_bits;
  assign regs_55_io_init = 64'h0;
  assign regs_55_io_enable = 1'h1;
  assign regs_55_clock = clock;
  assign regs_55_reset = reset;
  assign regs_56_io_in = io_argOuts_53_bits;
  assign regs_56_io_init = 64'h0;
  assign regs_56_io_enable = 1'h1;
  assign regs_56_clock = clock;
  assign regs_56_reset = reset;
  assign regs_57_io_in = io_argOuts_54_bits;
  assign regs_57_io_init = 64'h0;
  assign regs_57_io_enable = 1'h1;
  assign regs_57_clock = clock;
  assign regs_57_reset = reset;
  assign regs_58_io_in = io_argOuts_55_bits;
  assign regs_58_io_init = 64'h0;
  assign regs_58_io_enable = 1'h1;
  assign regs_58_clock = clock;
  assign regs_58_reset = reset;
  assign regs_59_io_in = io_argOuts_56_bits;
  assign regs_59_io_init = 64'h0;
  assign regs_59_io_enable = 1'h1;
  assign regs_59_clock = clock;
  assign regs_59_reset = reset;
  assign regs_60_io_in = io_argOuts_57_bits;
  assign regs_60_io_init = 64'h0;
  assign regs_60_io_enable = 1'h1;
  assign regs_60_clock = clock;
  assign regs_60_reset = reset;
  assign regs_61_io_in = io_argOuts_58_bits;
  assign regs_61_io_init = 64'h0;
  assign regs_61_io_enable = 1'h1;
  assign regs_61_clock = clock;
  assign regs_61_reset = reset;
  assign regs_62_io_in = io_argOuts_59_bits;
  assign regs_62_io_init = 64'h0;
  assign regs_62_io_enable = 1'h1;
  assign regs_62_clock = clock;
  assign regs_62_reset = reset;
  assign regs_63_io_in = io_argOuts_60_bits;
  assign regs_63_io_init = 64'h0;
  assign regs_63_io_enable = 1'h1;
  assign regs_63_clock = clock;
  assign regs_63_reset = reset;
  assign regs_64_io_in = io_argOuts_61_bits;
  assign regs_64_io_init = 64'h0;
  assign regs_64_io_enable = 1'h1;
  assign regs_64_clock = clock;
  assign regs_64_reset = reset;
  assign regs_65_io_in = io_argOuts_62_bits;
  assign regs_65_io_init = 64'h0;
  assign regs_65_io_enable = 1'h1;
  assign regs_65_clock = clock;
  assign regs_65_reset = reset;
  assign regs_66_io_in = io_argOuts_63_bits;
  assign regs_66_io_init = 64'h0;
  assign regs_66_io_enable = 1'h1;
  assign regs_66_clock = clock;
  assign regs_66_reset = reset;
  assign regs_67_io_in = io_argOuts_64_bits;
  assign regs_67_io_init = 64'h0;
  assign regs_67_io_enable = 1'h1;
  assign regs_67_clock = clock;
  assign regs_67_reset = reset;
  assign regs_68_io_in = io_argOuts_65_bits;
  assign regs_68_io_init = 64'h0;
  assign regs_68_io_enable = 1'h1;
  assign regs_68_clock = clock;
  assign regs_68_reset = reset;
  assign regs_69_io_in = io_argOuts_66_bits;
  assign regs_69_io_init = 64'h0;
  assign regs_69_io_enable = 1'h1;
  assign regs_69_clock = clock;
  assign regs_69_reset = reset;
  assign regs_70_io_in = io_argOuts_67_bits;
  assign regs_70_io_init = 64'h0;
  assign regs_70_io_enable = 1'h1;
  assign regs_70_clock = clock;
  assign regs_70_reset = reset;
  assign regs_71_io_in = io_argOuts_68_bits;
  assign regs_71_io_init = 64'h0;
  assign regs_71_io_enable = 1'h1;
  assign regs_71_clock = clock;
  assign regs_71_reset = reset;
  assign regs_72_io_in = io_argOuts_69_bits;
  assign regs_72_io_init = 64'h0;
  assign regs_72_io_enable = 1'h1;
  assign regs_72_clock = clock;
  assign regs_72_reset = reset;
  assign regs_73_io_in = io_argOuts_70_bits;
  assign regs_73_io_init = 64'h0;
  assign regs_73_io_enable = 1'h1;
  assign regs_73_clock = clock;
  assign regs_73_reset = reset;
  assign regs_74_io_in = io_argOuts_71_bits;
  assign regs_74_io_init = 64'h0;
  assign regs_74_io_enable = 1'h1;
  assign regs_74_clock = clock;
  assign regs_74_reset = reset;
  assign regs_75_io_in = io_argOuts_72_bits;
  assign regs_75_io_init = 64'h0;
  assign regs_75_io_enable = 1'h1;
  assign regs_75_clock = clock;
  assign regs_75_reset = reset;
  assign regs_76_io_in = io_argOuts_73_bits;
  assign regs_76_io_init = 64'h0;
  assign regs_76_io_enable = 1'h1;
  assign regs_76_clock = clock;
  assign regs_76_reset = reset;
  assign regs_77_io_in = io_argOuts_74_bits;
  assign regs_77_io_init = 64'h0;
  assign regs_77_io_enable = 1'h1;
  assign regs_77_clock = clock;
  assign regs_77_reset = reset;
  assign regs_78_io_in = io_argOuts_75_bits;
  assign regs_78_io_init = 64'h0;
  assign regs_78_io_enable = 1'h1;
  assign regs_78_clock = clock;
  assign regs_78_reset = reset;
  assign regs_79_io_in = io_argOuts_76_bits;
  assign regs_79_io_init = 64'h0;
  assign regs_79_io_enable = 1'h1;
  assign regs_79_clock = clock;
  assign regs_79_reset = reset;
  assign regs_80_io_in = io_argOuts_77_bits;
  assign regs_80_io_init = 64'h0;
  assign regs_80_io_enable = 1'h1;
  assign regs_80_clock = clock;
  assign regs_80_reset = reset;
  assign regs_81_io_in = io_argOuts_78_bits;
  assign regs_81_io_init = 64'h0;
  assign regs_81_io_enable = 1'h1;
  assign regs_81_clock = clock;
  assign regs_81_reset = reset;
  assign regs_82_io_in = io_argOuts_79_bits;
  assign regs_82_io_init = 64'h0;
  assign regs_82_io_enable = 1'h1;
  assign regs_82_clock = clock;
  assign regs_82_reset = reset;
  assign regs_83_io_in = io_argOuts_80_bits;
  assign regs_83_io_init = 64'h0;
  assign regs_83_io_enable = 1'h1;
  assign regs_83_clock = clock;
  assign regs_83_reset = reset;
  assign regs_84_io_in = io_argOuts_81_bits;
  assign regs_84_io_init = 64'h0;
  assign regs_84_io_enable = 1'h1;
  assign regs_84_clock = clock;
  assign regs_84_reset = reset;
  assign regs_85_io_in = io_argOuts_82_bits;
  assign regs_85_io_init = 64'h0;
  assign regs_85_io_enable = 1'h1;
  assign regs_85_clock = clock;
  assign regs_85_reset = reset;
  assign regs_86_io_in = io_argOuts_83_bits;
  assign regs_86_io_init = 64'h0;
  assign regs_86_io_enable = 1'h1;
  assign regs_86_clock = clock;
  assign regs_86_reset = reset;
  assign regs_87_io_in = io_argOuts_84_bits;
  assign regs_87_io_init = 64'h0;
  assign regs_87_io_enable = 1'h1;
  assign regs_87_clock = clock;
  assign regs_87_reset = reset;
  assign regs_88_io_in = io_argOuts_85_bits;
  assign regs_88_io_init = 64'h0;
  assign regs_88_io_enable = 1'h1;
  assign regs_88_clock = clock;
  assign regs_88_reset = reset;
  assign regs_89_io_in = io_argOuts_86_bits;
  assign regs_89_io_init = 64'h0;
  assign regs_89_io_enable = 1'h1;
  assign regs_89_clock = clock;
  assign regs_89_reset = reset;
  assign regs_90_io_in = io_argOuts_87_bits;
  assign regs_90_io_init = 64'h0;
  assign regs_90_io_enable = 1'h1;
  assign regs_90_clock = clock;
  assign regs_90_reset = reset;
  assign regs_91_io_in = io_argOuts_88_bits;
  assign regs_91_io_init = 64'h0;
  assign regs_91_io_enable = 1'h1;
  assign regs_91_clock = clock;
  assign regs_91_reset = reset;
  assign regs_92_io_in = io_argOuts_89_bits;
  assign regs_92_io_init = 64'h0;
  assign regs_92_io_enable = 1'h1;
  assign regs_92_clock = clock;
  assign regs_92_reset = reset;
  assign regs_93_io_in = io_argOuts_90_bits;
  assign regs_93_io_init = 64'h0;
  assign regs_93_io_enable = 1'h1;
  assign regs_93_clock = clock;
  assign regs_93_reset = reset;
  assign regs_94_io_in = io_argOuts_91_bits;
  assign regs_94_io_init = 64'h0;
  assign regs_94_io_enable = 1'h1;
  assign regs_94_clock = clock;
  assign regs_94_reset = reset;
  assign regs_95_io_in = io_argOuts_92_bits;
  assign regs_95_io_init = 64'h0;
  assign regs_95_io_enable = 1'h1;
  assign regs_95_clock = clock;
  assign regs_95_reset = reset;
  assign regs_96_io_in = io_argOuts_93_bits;
  assign regs_96_io_init = 64'h0;
  assign regs_96_io_enable = 1'h1;
  assign regs_96_clock = clock;
  assign regs_96_reset = reset;
  assign regs_97_io_in = io_argOuts_94_bits;
  assign regs_97_io_init = 64'h0;
  assign regs_97_io_enable = 1'h1;
  assign regs_97_clock = clock;
  assign regs_97_reset = reset;
  assign regs_98_io_in = io_argOuts_95_bits;
  assign regs_98_io_init = 64'h0;
  assign regs_98_io_enable = 1'h1;
  assign regs_98_clock = clock;
  assign regs_98_reset = reset;
  assign regs_99_io_in = io_argOuts_96_bits;
  assign regs_99_io_init = 64'h0;
  assign regs_99_io_enable = 1'h1;
  assign regs_99_clock = clock;
  assign regs_99_reset = reset;
  assign regs_100_io_in = io_argOuts_97_bits;
  assign regs_100_io_init = 64'h0;
  assign regs_100_io_enable = 1'h1;
  assign regs_100_clock = clock;
  assign regs_100_reset = reset;
  assign regs_101_io_in = io_argOuts_98_bits;
  assign regs_101_io_init = 64'h0;
  assign regs_101_io_enable = 1'h1;
  assign regs_101_clock = clock;
  assign regs_101_reset = reset;
  assign regs_102_io_in = io_argOuts_99_bits;
  assign regs_102_io_init = 64'h0;
  assign regs_102_io_enable = 1'h1;
  assign regs_102_clock = clock;
  assign regs_102_reset = reset;
  assign regs_103_io_in = io_argOuts_100_bits;
  assign regs_103_io_init = 64'h0;
  assign regs_103_io_enable = 1'h1;
  assign regs_103_clock = clock;
  assign regs_103_reset = reset;
  assign regs_104_io_in = io_argOuts_101_bits;
  assign regs_104_io_init = 64'h0;
  assign regs_104_io_enable = 1'h1;
  assign regs_104_clock = clock;
  assign regs_104_reset = reset;
  assign regs_105_io_in = io_argOuts_102_bits;
  assign regs_105_io_init = 64'h0;
  assign regs_105_io_enable = 1'h1;
  assign regs_105_clock = clock;
  assign regs_105_reset = reset;
  assign regs_106_io_in = io_argOuts_103_bits;
  assign regs_106_io_init = 64'h0;
  assign regs_106_io_enable = 1'h1;
  assign regs_106_clock = clock;
  assign regs_106_reset = reset;
  assign regs_107_io_in = io_argOuts_104_bits;
  assign regs_107_io_init = 64'h0;
  assign regs_107_io_enable = 1'h1;
  assign regs_107_clock = clock;
  assign regs_107_reset = reset;
  assign regs_108_io_in = io_argOuts_105_bits;
  assign regs_108_io_init = 64'h0;
  assign regs_108_io_enable = 1'h1;
  assign regs_108_clock = clock;
  assign regs_108_reset = reset;
  assign regs_109_io_in = io_argOuts_106_bits;
  assign regs_109_io_init = 64'h0;
  assign regs_109_io_enable = 1'h1;
  assign regs_109_clock = clock;
  assign regs_109_reset = reset;
  assign regs_110_io_in = io_argOuts_107_bits;
  assign regs_110_io_init = 64'h0;
  assign regs_110_io_enable = 1'h1;
  assign regs_110_clock = clock;
  assign regs_110_reset = reset;
  assign regs_111_io_in = io_argOuts_108_bits;
  assign regs_111_io_init = 64'h0;
  assign regs_111_io_enable = 1'h1;
  assign regs_111_clock = clock;
  assign regs_111_reset = reset;
  assign regs_112_io_in = io_argOuts_109_bits;
  assign regs_112_io_init = 64'h0;
  assign regs_112_io_enable = 1'h1;
  assign regs_112_clock = clock;
  assign regs_112_reset = reset;
  assign regs_113_io_in = io_argOuts_110_bits;
  assign regs_113_io_init = 64'h0;
  assign regs_113_io_enable = 1'h1;
  assign regs_113_clock = clock;
  assign regs_113_reset = reset;
  assign regs_114_io_in = io_argOuts_111_bits;
  assign regs_114_io_init = 64'h0;
  assign regs_114_io_enable = 1'h1;
  assign regs_114_clock = clock;
  assign regs_114_reset = reset;
  assign regs_115_io_in = io_argOuts_112_bits;
  assign regs_115_io_init = 64'h0;
  assign regs_115_io_enable = 1'h1;
  assign regs_115_clock = clock;
  assign regs_115_reset = reset;
  assign regs_116_io_in = io_argOuts_113_bits;
  assign regs_116_io_init = 64'h0;
  assign regs_116_io_enable = 1'h1;
  assign regs_116_clock = clock;
  assign regs_116_reset = reset;
  assign regs_117_io_in = io_argOuts_114_bits;
  assign regs_117_io_init = 64'h0;
  assign regs_117_io_enable = 1'h1;
  assign regs_117_clock = clock;
  assign regs_117_reset = reset;
  assign regs_118_io_in = io_argOuts_115_bits;
  assign regs_118_io_init = 64'h0;
  assign regs_118_io_enable = 1'h1;
  assign regs_118_clock = clock;
  assign regs_118_reset = reset;
  assign regs_119_io_in = 64'h0;
  assign regs_119_io_init = 64'h0;
  assign regs_119_io_enable = 1'h1;
  assign regs_119_clock = clock;
  assign regs_119_reset = reset;
  assign regs_120_io_in = 64'h0;
  assign regs_120_io_init = 64'h0;
  assign regs_120_io_enable = 1'h1;
  assign regs_120_clock = clock;
  assign regs_120_reset = reset;
  assign regs_121_io_in = 64'h0;
  assign regs_121_io_init = 64'h0;
  assign regs_121_io_enable = 1'h1;
  assign regs_121_clock = clock;
  assign regs_121_reset = reset;
  assign regs_122_io_in = 64'h0;
  assign regs_122_io_init = 64'h0;
  assign regs_122_io_enable = 1'h1;
  assign regs_122_clock = clock;
  assign regs_122_reset = reset;
  assign regs_123_io_in = 64'h0;
  assign regs_123_io_init = 64'h0;
  assign regs_123_io_enable = 1'h1;
  assign regs_123_clock = clock;
  assign regs_123_reset = reset;
  assign regs_124_io_in = 64'h0;
  assign regs_124_io_init = 64'h0;
  assign regs_124_io_enable = 1'h1;
  assign regs_124_clock = clock;
  assign regs_124_reset = reset;
  assign regs_125_io_in = 64'h0;
  assign regs_125_io_init = 64'h0;
  assign regs_125_io_enable = 1'h1;
  assign regs_125_clock = clock;
  assign regs_125_reset = reset;
  assign regs_126_io_in = 64'h0;
  assign regs_126_io_init = 64'h0;
  assign regs_126_io_enable = 1'h1;
  assign regs_126_clock = clock;
  assign regs_126_reset = reset;
  assign regs_127_io_in = 64'h0;
  assign regs_127_io_init = 64'h0;
  assign regs_127_io_enable = 1'h1;
  assign regs_127_clock = clock;
  assign regs_127_reset = reset;
  assign regs_128_io_in = 64'h0;
  assign regs_128_io_init = 64'h0;
  assign regs_128_io_enable = 1'h1;
  assign regs_128_clock = clock;
  assign regs_128_reset = reset;
  assign regs_129_io_in = 64'h0;
  assign regs_129_io_init = 64'h0;
  assign regs_129_io_enable = 1'h1;
  assign regs_129_clock = clock;
  assign regs_129_reset = reset;
  assign regs_130_io_in = 64'h0;
  assign regs_130_io_init = 64'h0;
  assign regs_130_io_enable = 1'h1;
  assign regs_130_clock = clock;
  assign regs_130_reset = reset;
  assign regs_131_io_in = 64'h0;
  assign regs_131_io_init = 64'h0;
  assign regs_131_io_enable = 1'h1;
  assign regs_131_clock = clock;
  assign regs_131_reset = reset;
  assign regs_132_io_in = 64'h0;
  assign regs_132_io_init = 64'h0;
  assign regs_132_io_enable = 1'h1;
  assign regs_132_clock = clock;
  assign regs_132_reset = reset;
  assign regs_133_io_in = 64'h0;
  assign regs_133_io_init = 64'h0;
  assign regs_133_io_enable = 1'h1;
  assign regs_133_clock = clock;
  assign regs_133_reset = reset;
  assign regs_134_io_in = 64'h0;
  assign regs_134_io_init = 64'h0;
  assign regs_134_io_enable = 1'h1;
  assign regs_134_clock = clock;
  assign regs_134_reset = reset;
  assign regs_135_io_in = 64'h0;
  assign regs_135_io_init = 64'h0;
  assign regs_135_io_enable = 1'h1;
  assign regs_135_clock = clock;
  assign regs_135_reset = reset;
  assign regs_136_io_in = 64'h0;
  assign regs_136_io_init = 64'h0;
  assign regs_136_io_enable = 1'h1;
  assign regs_136_clock = clock;
  assign regs_136_reset = reset;
  assign regs_137_io_in = 64'h0;
  assign regs_137_io_init = 64'h0;
  assign regs_137_io_enable = 1'h1;
  assign regs_137_clock = clock;
  assign regs_137_reset = reset;
  assign regs_138_io_in = 64'h0;
  assign regs_138_io_init = 64'h0;
  assign regs_138_io_enable = 1'h1;
  assign regs_138_clock = clock;
  assign regs_138_reset = reset;
  assign regs_139_io_in = 64'h0;
  assign regs_139_io_init = 64'h0;
  assign regs_139_io_enable = 1'h1;
  assign regs_139_clock = clock;
  assign regs_139_reset = reset;
  assign regs_140_io_in = 64'h0;
  assign regs_140_io_init = 64'h0;
  assign regs_140_io_enable = 1'h1;
  assign regs_140_clock = clock;
  assign regs_140_reset = reset;
  assign regs_141_io_in = 64'h0;
  assign regs_141_io_init = 64'h0;
  assign regs_141_io_enable = 1'h1;
  assign regs_141_clock = clock;
  assign regs_141_reset = reset;
  assign regs_142_io_in = 64'h0;
  assign regs_142_io_init = 64'h0;
  assign regs_142_io_enable = 1'h1;
  assign regs_142_clock = clock;
  assign regs_142_reset = reset;
  assign regs_143_io_in = 64'h0;
  assign regs_143_io_init = 64'h0;
  assign regs_143_io_enable = 1'h1;
  assign regs_143_clock = clock;
  assign regs_143_reset = reset;
  assign regs_144_io_in = 64'h0;
  assign regs_144_io_init = 64'h0;
  assign regs_144_io_enable = 1'h1;
  assign regs_144_clock = clock;
  assign regs_144_reset = reset;
  assign regs_145_io_in = 64'h0;
  assign regs_145_io_init = 64'h0;
  assign regs_145_io_enable = 1'h1;
  assign regs_145_clock = clock;
  assign regs_145_reset = reset;
  assign regs_146_io_in = 64'h0;
  assign regs_146_io_init = 64'h0;
  assign regs_146_io_enable = 1'h1;
  assign regs_146_clock = clock;
  assign regs_146_reset = reset;
  assign regs_147_io_in = 64'h0;
  assign regs_147_io_init = 64'h0;
  assign regs_147_io_enable = 1'h1;
  assign regs_147_clock = clock;
  assign regs_147_reset = reset;
  assign regs_148_io_in = 64'h0;
  assign regs_148_io_init = 64'h0;
  assign regs_148_io_enable = 1'h1;
  assign regs_148_clock = clock;
  assign regs_148_reset = reset;
  assign regs_149_io_in = 64'h0;
  assign regs_149_io_init = 64'h0;
  assign regs_149_io_enable = 1'h1;
  assign regs_149_clock = clock;
  assign regs_149_reset = reset;
  assign regs_150_io_in = 64'h0;
  assign regs_150_io_init = 64'h0;
  assign regs_150_io_enable = 1'h1;
  assign regs_150_clock = clock;
  assign regs_150_reset = reset;
  assign regs_151_io_in = 64'h0;
  assign regs_151_io_init = 64'h0;
  assign regs_151_io_enable = 1'h1;
  assign regs_151_clock = clock;
  assign regs_151_reset = reset;
  assign regs_152_io_in = 64'h0;
  assign regs_152_io_init = 64'h0;
  assign regs_152_io_enable = 1'h1;
  assign regs_152_clock = clock;
  assign regs_152_reset = reset;
  assign regs_153_io_in = 64'h0;
  assign regs_153_io_init = 64'h0;
  assign regs_153_io_enable = 1'h1;
  assign regs_153_clock = clock;
  assign regs_153_reset = reset;
  assign regs_154_io_in = 64'h0;
  assign regs_154_io_init = 64'h0;
  assign regs_154_io_enable = 1'h1;
  assign regs_154_clock = clock;
  assign regs_154_reset = reset;
  assign regs_155_io_in = 64'h0;
  assign regs_155_io_init = 64'h0;
  assign regs_155_io_enable = 1'h1;
  assign regs_155_clock = clock;
  assign regs_155_reset = reset;
  assign regs_156_io_in = 64'h0;
  assign regs_156_io_init = 64'h0;
  assign regs_156_io_enable = 1'h1;
  assign regs_156_clock = clock;
  assign regs_156_reset = reset;
  assign regs_157_io_in = 64'h0;
  assign regs_157_io_init = 64'h0;
  assign regs_157_io_enable = 1'h1;
  assign regs_157_clock = clock;
  assign regs_157_reset = reset;
  assign regs_158_io_in = 64'h0;
  assign regs_158_io_init = 64'h0;
  assign regs_158_io_enable = 1'h1;
  assign regs_158_clock = clock;
  assign regs_158_reset = reset;
  assign regs_159_io_in = 64'h0;
  assign regs_159_io_init = 64'h0;
  assign regs_159_io_enable = 1'h1;
  assign regs_159_clock = clock;
  assign regs_159_reset = reset;
  assign regs_160_io_in = 64'h0;
  assign regs_160_io_init = 64'h0;
  assign regs_160_io_enable = 1'h1;
  assign regs_160_clock = clock;
  assign regs_160_reset = reset;
  assign regs_161_io_in = 64'h0;
  assign regs_161_io_init = 64'h0;
  assign regs_161_io_enable = 1'h1;
  assign regs_161_clock = clock;
  assign regs_161_reset = reset;
  assign regs_162_io_in = 64'h0;
  assign regs_162_io_init = 64'h0;
  assign regs_162_io_enable = 1'h1;
  assign regs_162_clock = clock;
  assign regs_162_reset = reset;
  assign regs_163_io_in = 64'h0;
  assign regs_163_io_init = 64'h0;
  assign regs_163_io_enable = 1'h1;
  assign regs_163_clock = clock;
  assign regs_163_reset = reset;
  assign regs_164_io_in = 64'h0;
  assign regs_164_io_init = 64'h0;
  assign regs_164_io_enable = 1'h1;
  assign regs_164_clock = clock;
  assign regs_164_reset = reset;
  assign regs_165_io_in = 64'h0;
  assign regs_165_io_init = 64'h0;
  assign regs_165_io_enable = 1'h1;
  assign regs_165_clock = clock;
  assign regs_165_reset = reset;
  assign regs_166_io_in = 64'h0;
  assign regs_166_io_init = 64'h0;
  assign regs_166_io_enable = 1'h1;
  assign regs_166_clock = clock;
  assign regs_166_reset = reset;
  assign regs_167_io_in = 64'h0;
  assign regs_167_io_init = 64'h0;
  assign regs_167_io_enable = 1'h1;
  assign regs_167_clock = clock;
  assign regs_167_reset = reset;
  assign regs_168_io_in = 64'h0;
  assign regs_168_io_init = 64'h0;
  assign regs_168_io_enable = 1'h1;
  assign regs_168_clock = clock;
  assign regs_168_reset = reset;
  assign regs_169_io_in = 64'h0;
  assign regs_169_io_init = 64'h0;
  assign regs_169_io_enable = 1'h1;
  assign regs_169_clock = clock;
  assign regs_169_reset = reset;
  assign regs_170_io_in = 64'h0;
  assign regs_170_io_init = 64'h0;
  assign regs_170_io_enable = 1'h1;
  assign regs_170_clock = clock;
  assign regs_170_reset = reset;
  assign regs_171_io_in = 64'h0;
  assign regs_171_io_init = 64'h0;
  assign regs_171_io_enable = 1'h1;
  assign regs_171_clock = clock;
  assign regs_171_reset = reset;
  assign regs_172_io_in = 64'h0;
  assign regs_172_io_init = 64'h0;
  assign regs_172_io_enable = 1'h1;
  assign regs_172_clock = clock;
  assign regs_172_reset = reset;
  assign regs_173_io_in = 64'h0;
  assign regs_173_io_init = 64'h0;
  assign regs_173_io_enable = 1'h1;
  assign regs_173_clock = clock;
  assign regs_173_reset = reset;
  assign regs_174_io_in = 64'h0;
  assign regs_174_io_init = 64'h0;
  assign regs_174_io_enable = 1'h1;
  assign regs_174_clock = clock;
  assign regs_174_reset = reset;
  assign regs_175_io_in = 64'h0;
  assign regs_175_io_init = 64'h0;
  assign regs_175_io_enable = 1'h1;
  assign regs_175_clock = clock;
  assign regs_175_reset = reset;
  assign regs_176_io_in = 64'h0;
  assign regs_176_io_init = 64'h0;
  assign regs_176_io_enable = 1'h1;
  assign regs_176_clock = clock;
  assign regs_176_reset = reset;
  assign regs_177_io_in = 64'h0;
  assign regs_177_io_init = 64'h0;
  assign regs_177_io_enable = 1'h1;
  assign regs_177_clock = clock;
  assign regs_177_reset = reset;
  assign regs_178_io_in = 64'h0;
  assign regs_178_io_init = 64'h0;
  assign regs_178_io_enable = 1'h1;
  assign regs_178_clock = clock;
  assign regs_178_reset = reset;
  assign regs_179_io_in = 64'h0;
  assign regs_179_io_init = 64'h0;
  assign regs_179_io_enable = 1'h1;
  assign regs_179_clock = clock;
  assign regs_179_reset = reset;
  assign regs_180_io_in = 64'h0;
  assign regs_180_io_init = 64'h0;
  assign regs_180_io_enable = 1'h1;
  assign regs_180_clock = clock;
  assign regs_180_reset = reset;
  assign regs_181_io_in = 64'h0;
  assign regs_181_io_init = 64'h0;
  assign regs_181_io_enable = 1'h1;
  assign regs_181_clock = clock;
  assign regs_181_reset = reset;
  assign regs_182_io_in = 64'h0;
  assign regs_182_io_init = 64'h0;
  assign regs_182_io_enable = 1'h1;
  assign regs_182_clock = clock;
  assign regs_182_reset = reset;
  assign regs_183_io_in = 64'h0;
  assign regs_183_io_init = 64'h0;
  assign regs_183_io_enable = 1'h1;
  assign regs_183_clock = clock;
  assign regs_183_reset = reset;
  assign regs_184_io_in = 64'h0;
  assign regs_184_io_init = 64'h0;
  assign regs_184_io_enable = 1'h1;
  assign regs_184_clock = clock;
  assign regs_184_reset = reset;
  assign regs_185_io_in = 64'h0;
  assign regs_185_io_init = 64'h0;
  assign regs_185_io_enable = 1'h1;
  assign regs_185_clock = clock;
  assign regs_185_reset = reset;
  assign regs_186_io_in = 64'h0;
  assign regs_186_io_init = 64'h0;
  assign regs_186_io_enable = 1'h1;
  assign regs_186_clock = clock;
  assign regs_186_reset = reset;
  assign regs_187_io_in = 64'h0;
  assign regs_187_io_init = 64'h0;
  assign regs_187_io_enable = 1'h1;
  assign regs_187_clock = clock;
  assign regs_187_reset = reset;
  assign regs_188_io_in = 64'h0;
  assign regs_188_io_init = 64'h0;
  assign regs_188_io_enable = 1'h1;
  assign regs_188_clock = clock;
  assign regs_188_reset = reset;
  assign regs_189_io_in = 64'h0;
  assign regs_189_io_init = 64'h0;
  assign regs_189_io_enable = 1'h1;
  assign regs_189_clock = clock;
  assign regs_189_reset = reset;
  assign regs_190_io_in = 64'h0;
  assign regs_190_io_init = 64'h0;
  assign regs_190_io_enable = 1'h1;
  assign regs_190_clock = clock;
  assign regs_190_reset = reset;
  assign regs_191_io_in = 64'h0;
  assign regs_191_io_init = 64'h0;
  assign regs_191_io_enable = 1'h1;
  assign regs_191_clock = clock;
  assign regs_191_reset = reset;
  assign regs_192_io_in = 64'h0;
  assign regs_192_io_init = 64'h0;
  assign regs_192_io_enable = 1'h1;
  assign regs_192_clock = clock;
  assign regs_192_reset = reset;
  assign regs_193_io_in = 64'h0;
  assign regs_193_io_init = 64'h0;
  assign regs_193_io_enable = 1'h1;
  assign regs_193_clock = clock;
  assign regs_193_reset = reset;
  assign regs_194_io_in = 64'h0;
  assign regs_194_io_init = 64'h0;
  assign regs_194_io_enable = 1'h1;
  assign regs_194_clock = clock;
  assign regs_194_reset = reset;
  assign regs_195_io_in = 64'h0;
  assign regs_195_io_init = 64'h0;
  assign regs_195_io_enable = 1'h1;
  assign regs_195_clock = clock;
  assign regs_195_reset = reset;
  assign regs_196_io_in = 64'h0;
  assign regs_196_io_init = 64'h0;
  assign regs_196_io_enable = 1'h1;
  assign regs_196_clock = clock;
  assign regs_196_reset = reset;
  assign regs_197_io_in = 64'h0;
  assign regs_197_io_init = 64'h0;
  assign regs_197_io_enable = 1'h1;
  assign regs_197_clock = clock;
  assign regs_197_reset = reset;
  assign regs_198_io_in = 64'h0;
  assign regs_198_io_init = 64'h0;
  assign regs_198_io_enable = 1'h1;
  assign regs_198_clock = clock;
  assign regs_198_reset = reset;
  assign regs_199_io_in = 64'h0;
  assign regs_199_io_init = 64'h0;
  assign regs_199_io_enable = 1'h1;
  assign regs_199_clock = clock;
  assign regs_199_reset = reset;
  assign regs_200_io_in = 64'h0;
  assign regs_200_io_init = 64'h0;
  assign regs_200_io_enable = 1'h1;
  assign regs_200_clock = clock;
  assign regs_200_reset = reset;
  assign regs_201_io_in = 64'h0;
  assign regs_201_io_init = 64'h0;
  assign regs_201_io_enable = 1'h1;
  assign regs_201_clock = clock;
  assign regs_201_reset = reset;
  assign regs_202_io_in = 64'h0;
  assign regs_202_io_init = 64'h0;
  assign regs_202_io_enable = 1'h1;
  assign regs_202_clock = clock;
  assign regs_202_reset = reset;
  assign regs_203_io_in = 64'h0;
  assign regs_203_io_init = 64'h0;
  assign regs_203_io_enable = 1'h1;
  assign regs_203_clock = clock;
  assign regs_203_reset = reset;
  assign regs_204_io_in = 64'h0;
  assign regs_204_io_init = 64'h0;
  assign regs_204_io_enable = 1'h1;
  assign regs_204_clock = clock;
  assign regs_204_reset = reset;
  assign regs_205_io_in = 64'h0;
  assign regs_205_io_init = 64'h0;
  assign regs_205_io_enable = 1'h1;
  assign regs_205_clock = clock;
  assign regs_205_reset = reset;
  assign regs_206_io_in = 64'h0;
  assign regs_206_io_init = 64'h0;
  assign regs_206_io_enable = 1'h1;
  assign regs_206_clock = clock;
  assign regs_206_reset = reset;
  assign regs_207_io_in = 64'h0;
  assign regs_207_io_init = 64'h0;
  assign regs_207_io_enable = 1'h1;
  assign regs_207_clock = clock;
  assign regs_207_reset = reset;
  assign regs_208_io_in = 64'h0;
  assign regs_208_io_init = 64'h0;
  assign regs_208_io_enable = 1'h1;
  assign regs_208_clock = clock;
  assign regs_208_reset = reset;
  assign regs_209_io_in = 64'h0;
  assign regs_209_io_init = 64'h0;
  assign regs_209_io_enable = 1'h1;
  assign regs_209_clock = clock;
  assign regs_209_reset = reset;
  assign regs_210_io_in = 64'h0;
  assign regs_210_io_init = 64'h0;
  assign regs_210_io_enable = 1'h1;
  assign regs_210_clock = clock;
  assign regs_210_reset = reset;
  assign regs_211_io_in = 64'h0;
  assign regs_211_io_init = 64'h0;
  assign regs_211_io_enable = 1'h1;
  assign regs_211_clock = clock;
  assign regs_211_reset = reset;
  assign regs_212_io_in = 64'h0;
  assign regs_212_io_init = 64'h0;
  assign regs_212_io_enable = 1'h1;
  assign regs_212_clock = clock;
  assign regs_212_reset = reset;
  assign regs_213_io_in = 64'h0;
  assign regs_213_io_init = 64'h0;
  assign regs_213_io_enable = 1'h1;
  assign regs_213_clock = clock;
  assign regs_213_reset = reset;
  assign regs_214_io_in = 64'h0;
  assign regs_214_io_init = 64'h0;
  assign regs_214_io_enable = 1'h1;
  assign regs_214_clock = clock;
  assign regs_214_reset = reset;
  assign regs_215_io_in = 64'h0;
  assign regs_215_io_init = 64'h0;
  assign regs_215_io_enable = 1'h1;
  assign regs_215_clock = clock;
  assign regs_215_reset = reset;
  assign regs_216_io_in = 64'h0;
  assign regs_216_io_init = 64'h0;
  assign regs_216_io_enable = 1'h1;
  assign regs_216_clock = clock;
  assign regs_216_reset = reset;
  assign regs_217_io_in = 64'h0;
  assign regs_217_io_init = 64'h0;
  assign regs_217_io_enable = 1'h1;
  assign regs_217_clock = clock;
  assign regs_217_reset = reset;
  assign regs_218_io_in = 64'h0;
  assign regs_218_io_init = 64'h0;
  assign regs_218_io_enable = 1'h1;
  assign regs_218_clock = clock;
  assign regs_218_reset = reset;
  assign regs_219_io_in = 64'h0;
  assign regs_219_io_init = 64'h0;
  assign regs_219_io_enable = 1'h1;
  assign regs_219_clock = clock;
  assign regs_219_reset = reset;
  assign regs_220_io_in = 64'h0;
  assign regs_220_io_init = 64'h0;
  assign regs_220_io_enable = 1'h1;
  assign regs_220_clock = clock;
  assign regs_220_reset = reset;
  assign regs_221_io_in = 64'h0;
  assign regs_221_io_init = 64'h0;
  assign regs_221_io_enable = 1'h1;
  assign regs_221_clock = clock;
  assign regs_221_reset = reset;
  assign regs_222_io_in = 64'h0;
  assign regs_222_io_init = 64'h0;
  assign regs_222_io_enable = 1'h1;
  assign regs_222_clock = clock;
  assign regs_222_reset = reset;
  assign regs_223_io_in = 64'h0;
  assign regs_223_io_init = 64'h0;
  assign regs_223_io_enable = 1'h1;
  assign regs_223_clock = clock;
  assign regs_223_reset = reset;
  assign regs_224_io_in = 64'h0;
  assign regs_224_io_init = 64'h0;
  assign regs_224_io_enable = 1'h1;
  assign regs_224_clock = clock;
  assign regs_224_reset = reset;
  assign regs_225_io_in = 64'h0;
  assign regs_225_io_init = 64'h0;
  assign regs_225_io_enable = 1'h1;
  assign regs_225_clock = clock;
  assign regs_225_reset = reset;
  assign regs_226_io_in = 64'h0;
  assign regs_226_io_init = 64'h0;
  assign regs_226_io_enable = 1'h1;
  assign regs_226_clock = clock;
  assign regs_226_reset = reset;
  assign regs_227_io_in = 64'h0;
  assign regs_227_io_init = 64'h0;
  assign regs_227_io_enable = 1'h1;
  assign regs_227_clock = clock;
  assign regs_227_reset = reset;
  assign regs_228_io_in = 64'h0;
  assign regs_228_io_init = 64'h0;
  assign regs_228_io_enable = 1'h1;
  assign regs_228_clock = clock;
  assign regs_228_reset = reset;
  assign regs_229_io_in = 64'h0;
  assign regs_229_io_init = 64'h0;
  assign regs_229_io_enable = 1'h1;
  assign regs_229_clock = clock;
  assign regs_229_reset = reset;
  assign regs_230_io_in = 64'h0;
  assign regs_230_io_init = 64'h0;
  assign regs_230_io_enable = 1'h1;
  assign regs_230_clock = clock;
  assign regs_230_reset = reset;
  assign regs_231_io_in = 64'h0;
  assign regs_231_io_init = 64'h0;
  assign regs_231_io_enable = 1'h1;
  assign regs_231_clock = clock;
  assign regs_231_reset = reset;
  assign regs_232_io_in = 64'h0;
  assign regs_232_io_init = 64'h0;
  assign regs_232_io_enable = 1'h1;
  assign regs_232_clock = clock;
  assign regs_232_reset = reset;
  assign regs_233_io_in = 64'h0;
  assign regs_233_io_init = 64'h0;
  assign regs_233_io_enable = 1'h1;
  assign regs_233_clock = clock;
  assign regs_233_reset = reset;
  assign regs_234_io_in = 64'h0;
  assign regs_234_io_init = 64'h0;
  assign regs_234_io_enable = 1'h1;
  assign regs_234_clock = clock;
  assign regs_234_reset = reset;
  assign regs_235_io_in = 64'h0;
  assign regs_235_io_init = 64'h0;
  assign regs_235_io_enable = 1'h1;
  assign regs_235_clock = clock;
  assign regs_235_reset = reset;
  assign regs_236_io_in = 64'h0;
  assign regs_236_io_init = 64'h0;
  assign regs_236_io_enable = 1'h1;
  assign regs_236_clock = clock;
  assign regs_236_reset = reset;
  assign regs_237_io_in = 64'h0;
  assign regs_237_io_init = 64'h0;
  assign regs_237_io_enable = 1'h1;
  assign regs_237_clock = clock;
  assign regs_237_reset = reset;
  assign regs_238_io_in = 64'h0;
  assign regs_238_io_init = 64'h0;
  assign regs_238_io_enable = 1'h1;
  assign regs_238_clock = clock;
  assign regs_238_reset = reset;
  assign regs_239_io_in = 64'h0;
  assign regs_239_io_init = 64'h0;
  assign regs_239_io_enable = 1'h1;
  assign regs_239_clock = clock;
  assign regs_239_reset = reset;
  assign regs_240_io_in = 64'h0;
  assign regs_240_io_init = 64'h0;
  assign regs_240_io_enable = 1'h1;
  assign regs_240_clock = clock;
  assign regs_240_reset = reset;
  assign regs_241_io_in = 64'h0;
  assign regs_241_io_init = 64'h0;
  assign regs_241_io_enable = 1'h1;
  assign regs_241_clock = clock;
  assign regs_241_reset = reset;
  assign regs_242_io_in = 64'h0;
  assign regs_242_io_init = 64'h0;
  assign regs_242_io_enable = 1'h1;
  assign regs_242_clock = clock;
  assign regs_242_reset = reset;
  assign regs_243_io_in = 64'h0;
  assign regs_243_io_init = 64'h0;
  assign regs_243_io_enable = 1'h1;
  assign regs_243_clock = clock;
  assign regs_243_reset = reset;
  assign regs_244_io_in = 64'h0;
  assign regs_244_io_init = 64'h0;
  assign regs_244_io_enable = 1'h1;
  assign regs_244_clock = clock;
  assign regs_244_reset = reset;
  assign regs_245_io_in = 64'h0;
  assign regs_245_io_init = 64'h0;
  assign regs_245_io_enable = 1'h1;
  assign regs_245_clock = clock;
  assign regs_245_reset = reset;
  assign regs_246_io_in = 64'h0;
  assign regs_246_io_init = 64'h0;
  assign regs_246_io_enable = 1'h1;
  assign regs_246_clock = clock;
  assign regs_246_reset = reset;
  assign regs_247_io_in = 64'h0;
  assign regs_247_io_init = 64'h0;
  assign regs_247_io_enable = 1'h1;
  assign regs_247_clock = clock;
  assign regs_247_reset = reset;
  assign regs_248_io_in = 64'h0;
  assign regs_248_io_init = 64'h0;
  assign regs_248_io_enable = 1'h1;
  assign regs_248_clock = clock;
  assign regs_248_reset = reset;
  assign regs_249_io_in = 64'h0;
  assign regs_249_io_init = 64'h0;
  assign regs_249_io_enable = 1'h1;
  assign regs_249_clock = clock;
  assign regs_249_reset = reset;
  assign regs_250_io_in = 64'h0;
  assign regs_250_io_init = 64'h0;
  assign regs_250_io_enable = 1'h1;
  assign regs_250_clock = clock;
  assign regs_250_reset = reset;
  assign regs_251_io_in = 64'h0;
  assign regs_251_io_init = 64'h0;
  assign regs_251_io_enable = 1'h1;
  assign regs_251_clock = clock;
  assign regs_251_reset = reset;
  assign regs_252_io_in = 64'h0;
  assign regs_252_io_init = 64'h0;
  assign regs_252_io_enable = 1'h1;
  assign regs_252_clock = clock;
  assign regs_252_reset = reset;
  assign regs_253_io_in = 64'h0;
  assign regs_253_io_init = 64'h0;
  assign regs_253_io_enable = 1'h1;
  assign regs_253_clock = clock;
  assign regs_253_reset = reset;
  assign regs_254_io_in = 64'h0;
  assign regs_254_io_init = 64'h0;
  assign regs_254_io_enable = 1'h1;
  assign regs_254_clock = clock;
  assign regs_254_reset = reset;
  assign regs_255_io_in = 64'h0;
  assign regs_255_io_init = 64'h0;
  assign regs_255_io_enable = 1'h1;
  assign regs_255_clock = clock;
  assign regs_255_reset = reset;
  assign regs_256_io_in = 64'h0;
  assign regs_256_io_init = 64'h0;
  assign regs_256_io_enable = 1'h1;
  assign regs_256_clock = clock;
  assign regs_256_reset = reset;
  assign regs_257_io_in = 64'h0;
  assign regs_257_io_init = 64'h0;
  assign regs_257_io_enable = 1'h1;
  assign regs_257_clock = clock;
  assign regs_257_reset = reset;
  assign regs_258_io_in = 64'h0;
  assign regs_258_io_init = 64'h0;
  assign regs_258_io_enable = 1'h1;
  assign regs_258_clock = clock;
  assign regs_258_reset = reset;
  assign regs_259_io_in = 64'h0;
  assign regs_259_io_init = 64'h0;
  assign regs_259_io_enable = 1'h1;
  assign regs_259_clock = clock;
  assign regs_259_reset = reset;
  assign regs_260_io_in = 64'h0;
  assign regs_260_io_init = 64'h0;
  assign regs_260_io_enable = 1'h1;
  assign regs_260_clock = clock;
  assign regs_260_reset = reset;
  assign regs_261_io_in = 64'h0;
  assign regs_261_io_init = 64'h0;
  assign regs_261_io_enable = 1'h1;
  assign regs_261_clock = clock;
  assign regs_261_reset = reset;
  assign regs_262_io_in = 64'h0;
  assign regs_262_io_init = 64'h0;
  assign regs_262_io_enable = 1'h1;
  assign regs_262_clock = clock;
  assign regs_262_reset = reset;
  assign regs_263_io_in = 64'h0;
  assign regs_263_io_init = 64'h0;
  assign regs_263_io_enable = 1'h1;
  assign regs_263_clock = clock;
  assign regs_263_reset = reset;
  assign regs_264_io_in = 64'h0;
  assign regs_264_io_init = 64'h0;
  assign regs_264_io_enable = 1'h1;
  assign regs_264_clock = clock;
  assign regs_264_reset = reset;
  assign regs_265_io_in = 64'h0;
  assign regs_265_io_init = 64'h0;
  assign regs_265_io_enable = 1'h1;
  assign regs_265_clock = clock;
  assign regs_265_reset = reset;
  assign regs_266_io_in = 64'h0;
  assign regs_266_io_init = 64'h0;
  assign regs_266_io_enable = 1'h1;
  assign regs_266_clock = clock;
  assign regs_266_reset = reset;
  assign regs_267_io_in = 64'h0;
  assign regs_267_io_init = 64'h0;
  assign regs_267_io_enable = 1'h1;
  assign regs_267_clock = clock;
  assign regs_267_reset = reset;
  assign regs_268_io_in = 64'h0;
  assign regs_268_io_init = 64'h0;
  assign regs_268_io_enable = 1'h1;
  assign regs_268_clock = clock;
  assign regs_268_reset = reset;
  assign regs_269_io_in = 64'h0;
  assign regs_269_io_init = 64'h0;
  assign regs_269_io_enable = 1'h1;
  assign regs_269_clock = clock;
  assign regs_269_reset = reset;
  assign regs_270_io_in = 64'h0;
  assign regs_270_io_init = 64'h0;
  assign regs_270_io_enable = 1'h1;
  assign regs_270_clock = clock;
  assign regs_270_reset = reset;
  assign regs_271_io_in = 64'h0;
  assign regs_271_io_init = 64'h0;
  assign regs_271_io_enable = 1'h1;
  assign regs_271_clock = clock;
  assign regs_271_reset = reset;
  assign regs_272_io_in = 64'h0;
  assign regs_272_io_init = 64'h0;
  assign regs_272_io_enable = 1'h1;
  assign regs_272_clock = clock;
  assign regs_272_reset = reset;
  assign regs_273_io_in = 64'h0;
  assign regs_273_io_init = 64'h0;
  assign regs_273_io_enable = 1'h1;
  assign regs_273_clock = clock;
  assign regs_273_reset = reset;
  assign regs_274_io_in = 64'h0;
  assign regs_274_io_init = 64'h0;
  assign regs_274_io_enable = 1'h1;
  assign regs_274_clock = clock;
  assign regs_274_reset = reset;
  assign regs_275_io_in = 64'h0;
  assign regs_275_io_init = 64'h0;
  assign regs_275_io_enable = 1'h1;
  assign regs_275_clock = clock;
  assign regs_275_reset = reset;
  assign regs_276_io_in = 64'h0;
  assign regs_276_io_init = 64'h0;
  assign regs_276_io_enable = 1'h1;
  assign regs_276_clock = clock;
  assign regs_276_reset = reset;
  assign regs_277_io_in = 64'h0;
  assign regs_277_io_init = 64'h0;
  assign regs_277_io_enable = 1'h1;
  assign regs_277_clock = clock;
  assign regs_277_reset = reset;
  assign regs_278_io_in = 64'h0;
  assign regs_278_io_init = 64'h0;
  assign regs_278_io_enable = 1'h1;
  assign regs_278_clock = clock;
  assign regs_278_reset = reset;
  assign regs_279_io_in = 64'h0;
  assign regs_279_io_init = 64'h0;
  assign regs_279_io_enable = 1'h1;
  assign regs_279_clock = clock;
  assign regs_279_reset = reset;
  assign regs_280_io_in = 64'h0;
  assign regs_280_io_init = 64'h0;
  assign regs_280_io_enable = 1'h1;
  assign regs_280_clock = clock;
  assign regs_280_reset = reset;
  assign regs_281_io_in = 64'h0;
  assign regs_281_io_init = 64'h0;
  assign regs_281_io_enable = 1'h1;
  assign regs_281_clock = clock;
  assign regs_281_reset = reset;
  assign regs_282_io_in = 64'h0;
  assign regs_282_io_init = 64'h0;
  assign regs_282_io_enable = 1'h1;
  assign regs_282_clock = clock;
  assign regs_282_reset = reset;
  assign regs_283_io_in = 64'h0;
  assign regs_283_io_init = 64'h0;
  assign regs_283_io_enable = 1'h1;
  assign regs_283_clock = clock;
  assign regs_283_reset = reset;
  assign regs_284_io_in = 64'h0;
  assign regs_284_io_init = 64'h0;
  assign regs_284_io_enable = 1'h1;
  assign regs_284_clock = clock;
  assign regs_284_reset = reset;
  assign regs_285_io_in = 64'h0;
  assign regs_285_io_init = 64'h0;
  assign regs_285_io_enable = 1'h1;
  assign regs_285_clock = clock;
  assign regs_285_reset = reset;
  assign regs_286_io_in = 64'h0;
  assign regs_286_io_init = 64'h0;
  assign regs_286_io_enable = 1'h1;
  assign regs_286_clock = clock;
  assign regs_286_reset = reset;
  assign regs_287_io_in = 64'h0;
  assign regs_287_io_init = 64'h0;
  assign regs_287_io_enable = 1'h1;
  assign regs_287_clock = clock;
  assign regs_287_reset = reset;
  assign regs_288_io_in = 64'h0;
  assign regs_288_io_init = 64'h0;
  assign regs_288_io_enable = 1'h1;
  assign regs_288_clock = clock;
  assign regs_288_reset = reset;
  assign regs_289_io_in = 64'h0;
  assign regs_289_io_init = 64'h0;
  assign regs_289_io_enable = 1'h1;
  assign regs_289_clock = clock;
  assign regs_289_reset = reset;
  assign regs_290_io_in = 64'h0;
  assign regs_290_io_init = 64'h0;
  assign regs_290_io_enable = 1'h1;
  assign regs_290_clock = clock;
  assign regs_290_reset = reset;
  assign regs_291_io_in = 64'h0;
  assign regs_291_io_init = 64'h0;
  assign regs_291_io_enable = 1'h1;
  assign regs_291_clock = clock;
  assign regs_291_reset = reset;
  assign regs_292_io_in = 64'h0;
  assign regs_292_io_init = 64'h0;
  assign regs_292_io_enable = 1'h1;
  assign regs_292_clock = clock;
  assign regs_292_reset = reset;
  assign regs_293_io_in = 64'h0;
  assign regs_293_io_init = 64'h0;
  assign regs_293_io_enable = 1'h1;
  assign regs_293_clock = clock;
  assign regs_293_reset = reset;
  assign regs_294_io_in = 64'h0;
  assign regs_294_io_init = 64'h0;
  assign regs_294_io_enable = 1'h1;
  assign regs_294_clock = clock;
  assign regs_294_reset = reset;
  assign regs_295_io_in = 64'h0;
  assign regs_295_io_init = 64'h0;
  assign regs_295_io_enable = 1'h1;
  assign regs_295_clock = clock;
  assign regs_295_reset = reset;
  assign regs_296_io_in = 64'h0;
  assign regs_296_io_init = 64'h0;
  assign regs_296_io_enable = 1'h1;
  assign regs_296_clock = clock;
  assign regs_296_reset = reset;
  assign regs_297_io_in = 64'h0;
  assign regs_297_io_init = 64'h0;
  assign regs_297_io_enable = 1'h1;
  assign regs_297_clock = clock;
  assign regs_297_reset = reset;
  assign regs_298_io_in = 64'h0;
  assign regs_298_io_init = 64'h0;
  assign regs_298_io_enable = 1'h1;
  assign regs_298_clock = clock;
  assign regs_298_reset = reset;
  assign regs_299_io_in = 64'h0;
  assign regs_299_io_init = 64'h0;
  assign regs_299_io_enable = 1'h1;
  assign regs_299_clock = clock;
  assign regs_299_reset = reset;
  assign regs_300_io_in = 64'h0;
  assign regs_300_io_init = 64'h0;
  assign regs_300_io_enable = 1'h1;
  assign regs_300_clock = clock;
  assign regs_300_reset = reset;
  assign regs_301_io_in = 64'h0;
  assign regs_301_io_init = 64'h0;
  assign regs_301_io_enable = 1'h1;
  assign regs_301_clock = clock;
  assign regs_301_reset = reset;
  assign regs_302_io_in = 64'h0;
  assign regs_302_io_init = 64'h0;
  assign regs_302_io_enable = 1'h1;
  assign regs_302_clock = clock;
  assign regs_302_reset = reset;
  assign regs_303_io_in = 64'h0;
  assign regs_303_io_init = 64'h0;
  assign regs_303_io_enable = 1'h1;
  assign regs_303_clock = clock;
  assign regs_303_reset = reset;
  assign regs_304_io_in = 64'h0;
  assign regs_304_io_init = 64'h0;
  assign regs_304_io_enable = 1'h1;
  assign regs_304_clock = clock;
  assign regs_304_reset = reset;
  assign regs_305_io_in = 64'h0;
  assign regs_305_io_init = 64'h0;
  assign regs_305_io_enable = 1'h1;
  assign regs_305_clock = clock;
  assign regs_305_reset = reset;
  assign regs_306_io_in = 64'h0;
  assign regs_306_io_init = 64'h0;
  assign regs_306_io_enable = 1'h1;
  assign regs_306_clock = clock;
  assign regs_306_reset = reset;
  assign regs_307_io_in = 64'h0;
  assign regs_307_io_init = 64'h0;
  assign regs_307_io_enable = 1'h1;
  assign regs_307_clock = clock;
  assign regs_307_reset = reset;
  assign regs_308_io_in = 64'h0;
  assign regs_308_io_init = 64'h0;
  assign regs_308_io_enable = 1'h1;
  assign regs_308_clock = clock;
  assign regs_308_reset = reset;
  assign regs_309_io_in = 64'h0;
  assign regs_309_io_init = 64'h0;
  assign regs_309_io_enable = 1'h1;
  assign regs_309_clock = clock;
  assign regs_309_reset = reset;
  assign regs_310_io_in = 64'h0;
  assign regs_310_io_init = 64'h0;
  assign regs_310_io_enable = 1'h1;
  assign regs_310_clock = clock;
  assign regs_310_reset = reset;
  assign regs_311_io_in = 64'h0;
  assign regs_311_io_init = 64'h0;
  assign regs_311_io_enable = 1'h1;
  assign regs_311_clock = clock;
  assign regs_311_reset = reset;
  assign regs_312_io_in = 64'h0;
  assign regs_312_io_init = 64'h0;
  assign regs_312_io_enable = 1'h1;
  assign regs_312_clock = clock;
  assign regs_312_reset = reset;
  assign regs_313_io_in = 64'h0;
  assign regs_313_io_init = 64'h0;
  assign regs_313_io_enable = 1'h1;
  assign regs_313_clock = clock;
  assign regs_313_reset = reset;
  assign regs_314_io_in = 64'h0;
  assign regs_314_io_init = 64'h0;
  assign regs_314_io_enable = 1'h1;
  assign regs_314_clock = clock;
  assign regs_314_reset = reset;
  assign regs_315_io_in = 64'h0;
  assign regs_315_io_init = 64'h0;
  assign regs_315_io_enable = 1'h1;
  assign regs_315_clock = clock;
  assign regs_315_reset = reset;
  assign regs_316_io_in = 64'h0;
  assign regs_316_io_init = 64'h0;
  assign regs_316_io_enable = 1'h1;
  assign regs_316_clock = clock;
  assign regs_316_reset = reset;
  assign regs_317_io_in = 64'h0;
  assign regs_317_io_init = 64'h0;
  assign regs_317_io_enable = 1'h1;
  assign regs_317_clock = clock;
  assign regs_317_reset = reset;
  assign regs_318_io_in = 64'h0;
  assign regs_318_io_init = 64'h0;
  assign regs_318_io_enable = 1'h1;
  assign regs_318_clock = clock;
  assign regs_318_reset = reset;
  assign regs_319_io_in = 64'h0;
  assign regs_319_io_init = 64'h0;
  assign regs_319_io_enable = 1'h1;
  assign regs_319_clock = clock;
  assign regs_319_reset = reset;
  assign regs_320_io_in = 64'h0;
  assign regs_320_io_init = 64'h0;
  assign regs_320_io_enable = 1'h1;
  assign regs_320_clock = clock;
  assign regs_320_reset = reset;
  assign regs_321_io_in = 64'h0;
  assign regs_321_io_init = 64'h0;
  assign regs_321_io_enable = 1'h1;
  assign regs_321_clock = clock;
  assign regs_321_reset = reset;
  assign regs_322_io_in = 64'h0;
  assign regs_322_io_init = 64'h0;
  assign regs_322_io_enable = 1'h1;
  assign regs_322_clock = clock;
  assign regs_322_reset = reset;
  assign regs_323_io_in = 64'h0;
  assign regs_323_io_init = 64'h0;
  assign regs_323_io_enable = 1'h1;
  assign regs_323_clock = clock;
  assign regs_323_reset = reset;
  assign regs_324_io_in = 64'h0;
  assign regs_324_io_init = 64'h0;
  assign regs_324_io_enable = 1'h1;
  assign regs_324_clock = clock;
  assign regs_324_reset = reset;
  assign regs_325_io_in = 64'h0;
  assign regs_325_io_init = 64'h0;
  assign regs_325_io_enable = 1'h1;
  assign regs_325_clock = clock;
  assign regs_325_reset = reset;
  assign regs_326_io_in = 64'h0;
  assign regs_326_io_init = 64'h0;
  assign regs_326_io_enable = 1'h1;
  assign regs_326_clock = clock;
  assign regs_326_reset = reset;
  assign regs_327_io_in = 64'h0;
  assign regs_327_io_init = 64'h0;
  assign regs_327_io_enable = 1'h1;
  assign regs_327_clock = clock;
  assign regs_327_reset = reset;
  assign regs_328_io_in = 64'h0;
  assign regs_328_io_init = 64'h0;
  assign regs_328_io_enable = 1'h1;
  assign regs_328_clock = clock;
  assign regs_328_reset = reset;
  assign regs_329_io_in = 64'h0;
  assign regs_329_io_init = 64'h0;
  assign regs_329_io_enable = 1'h1;
  assign regs_329_clock = clock;
  assign regs_329_reset = reset;
  assign regs_330_io_in = 64'h0;
  assign regs_330_io_init = 64'h0;
  assign regs_330_io_enable = 1'h1;
  assign regs_330_clock = clock;
  assign regs_330_reset = reset;
  assign regs_331_io_in = 64'h0;
  assign regs_331_io_init = 64'h0;
  assign regs_331_io_enable = 1'h1;
  assign regs_331_clock = clock;
  assign regs_331_reset = reset;
  assign regs_332_io_in = 64'h0;
  assign regs_332_io_init = 64'h0;
  assign regs_332_io_enable = 1'h1;
  assign regs_332_clock = clock;
  assign regs_332_reset = reset;
  assign regs_333_io_in = 64'h0;
  assign regs_333_io_init = 64'h0;
  assign regs_333_io_enable = 1'h1;
  assign regs_333_clock = clock;
  assign regs_333_reset = reset;
  assign regs_334_io_in = 64'h0;
  assign regs_334_io_init = 64'h0;
  assign regs_334_io_enable = 1'h1;
  assign regs_334_clock = clock;
  assign regs_334_reset = reset;
  assign regs_335_io_in = 64'h0;
  assign regs_335_io_init = 64'h0;
  assign regs_335_io_enable = 1'h1;
  assign regs_335_clock = clock;
  assign regs_335_reset = reset;
  assign regs_336_io_in = 64'h0;
  assign regs_336_io_init = 64'h0;
  assign regs_336_io_enable = 1'h1;
  assign regs_336_clock = clock;
  assign regs_336_reset = reset;
  assign regs_337_io_in = 64'h0;
  assign regs_337_io_init = 64'h0;
  assign regs_337_io_enable = 1'h1;
  assign regs_337_clock = clock;
  assign regs_337_reset = reset;
  assign regs_338_io_in = 64'h0;
  assign regs_338_io_init = 64'h0;
  assign regs_338_io_enable = 1'h1;
  assign regs_338_clock = clock;
  assign regs_338_reset = reset;
  assign regs_339_io_in = 64'h0;
  assign regs_339_io_init = 64'h0;
  assign regs_339_io_enable = 1'h1;
  assign regs_339_clock = clock;
  assign regs_339_reset = reset;
  assign regs_340_io_in = 64'h0;
  assign regs_340_io_init = 64'h0;
  assign regs_340_io_enable = 1'h1;
  assign regs_340_clock = clock;
  assign regs_340_reset = reset;
  assign regs_341_io_in = 64'h0;
  assign regs_341_io_init = 64'h0;
  assign regs_341_io_enable = 1'h1;
  assign regs_341_clock = clock;
  assign regs_341_reset = reset;
  assign regs_342_io_in = 64'h0;
  assign regs_342_io_init = 64'h0;
  assign regs_342_io_enable = 1'h1;
  assign regs_342_clock = clock;
  assign regs_342_reset = reset;
  assign regs_343_io_in = 64'h0;
  assign regs_343_io_init = 64'h0;
  assign regs_343_io_enable = 1'h1;
  assign regs_343_clock = clock;
  assign regs_343_reset = reset;
  assign regs_344_io_in = 64'h0;
  assign regs_344_io_init = 64'h0;
  assign regs_344_io_enable = 1'h1;
  assign regs_344_clock = clock;
  assign regs_344_reset = reset;
  assign regs_345_io_in = 64'h0;
  assign regs_345_io_init = 64'h0;
  assign regs_345_io_enable = 1'h1;
  assign regs_345_clock = clock;
  assign regs_345_reset = reset;
  assign regs_346_io_in = 64'h0;
  assign regs_346_io_init = 64'h0;
  assign regs_346_io_enable = 1'h1;
  assign regs_346_clock = clock;
  assign regs_346_reset = reset;
  assign regs_347_io_in = 64'h0;
  assign regs_347_io_init = 64'h0;
  assign regs_347_io_enable = 1'h1;
  assign regs_347_clock = clock;
  assign regs_347_reset = reset;
  assign regs_348_io_in = 64'h0;
  assign regs_348_io_init = 64'h0;
  assign regs_348_io_enable = 1'h1;
  assign regs_348_clock = clock;
  assign regs_348_reset = reset;
  assign regs_349_io_in = 64'h0;
  assign regs_349_io_init = 64'h0;
  assign regs_349_io_enable = 1'h1;
  assign regs_349_clock = clock;
  assign regs_349_reset = reset;
  assign regs_350_io_in = 64'h0;
  assign regs_350_io_init = 64'h0;
  assign regs_350_io_enable = 1'h1;
  assign regs_350_clock = clock;
  assign regs_350_reset = reset;
  assign regs_351_io_in = 64'h0;
  assign regs_351_io_init = 64'h0;
  assign regs_351_io_enable = 1'h1;
  assign regs_351_clock = clock;
  assign regs_351_reset = reset;
  assign regs_352_io_in = 64'h0;
  assign regs_352_io_init = 64'h0;
  assign regs_352_io_enable = 1'h1;
  assign regs_352_clock = clock;
  assign regs_352_reset = reset;
  assign regs_353_io_in = 64'h0;
  assign regs_353_io_init = 64'h0;
  assign regs_353_io_enable = 1'h1;
  assign regs_353_clock = clock;
  assign regs_353_reset = reset;
  assign regs_354_io_in = 64'h0;
  assign regs_354_io_init = 64'h0;
  assign regs_354_io_enable = 1'h1;
  assign regs_354_clock = clock;
  assign regs_354_reset = reset;
  assign regs_355_io_in = 64'h0;
  assign regs_355_io_init = 64'h0;
  assign regs_355_io_enable = 1'h1;
  assign regs_355_clock = clock;
  assign regs_355_reset = reset;
  assign regs_356_io_in = 64'h0;
  assign regs_356_io_init = 64'h0;
  assign regs_356_io_enable = 1'h1;
  assign regs_356_clock = clock;
  assign regs_356_reset = reset;
  assign regs_357_io_in = 64'h0;
  assign regs_357_io_init = 64'h0;
  assign regs_357_io_enable = 1'h1;
  assign regs_357_clock = clock;
  assign regs_357_reset = reset;
  assign regs_358_io_in = 64'h0;
  assign regs_358_io_init = 64'h0;
  assign regs_358_io_enable = 1'h1;
  assign regs_358_clock = clock;
  assign regs_358_reset = reset;
  assign regs_359_io_in = 64'h0;
  assign regs_359_io_init = 64'h0;
  assign regs_359_io_enable = 1'h1;
  assign regs_359_clock = clock;
  assign regs_359_reset = reset;
  assign regs_360_io_in = 64'h0;
  assign regs_360_io_init = 64'h0;
  assign regs_360_io_enable = 1'h1;
  assign regs_360_clock = clock;
  assign regs_360_reset = reset;
  assign regs_361_io_in = 64'h0;
  assign regs_361_io_init = 64'h0;
  assign regs_361_io_enable = 1'h1;
  assign regs_361_clock = clock;
  assign regs_361_reset = reset;
  assign regs_362_io_in = 64'h0;
  assign regs_362_io_init = 64'h0;
  assign regs_362_io_enable = 1'h1;
  assign regs_362_clock = clock;
  assign regs_362_reset = reset;
  assign regs_363_io_in = 64'h0;
  assign regs_363_io_init = 64'h0;
  assign regs_363_io_enable = 1'h1;
  assign regs_363_clock = clock;
  assign regs_363_reset = reset;
  assign regs_364_io_in = 64'h0;
  assign regs_364_io_init = 64'h0;
  assign regs_364_io_enable = 1'h1;
  assign regs_364_clock = clock;
  assign regs_364_reset = reset;
  assign regs_365_io_in = 64'h0;
  assign regs_365_io_init = 64'h0;
  assign regs_365_io_enable = 1'h1;
  assign regs_365_clock = clock;
  assign regs_365_reset = reset;
  assign regs_366_io_in = 64'h0;
  assign regs_366_io_init = 64'h0;
  assign regs_366_io_enable = 1'h1;
  assign regs_366_clock = clock;
  assign regs_366_reset = reset;
  assign regs_367_io_in = 64'h0;
  assign regs_367_io_init = 64'h0;
  assign regs_367_io_enable = 1'h1;
  assign regs_367_clock = clock;
  assign regs_367_reset = reset;
  assign regs_368_io_in = 64'h0;
  assign regs_368_io_init = 64'h0;
  assign regs_368_io_enable = 1'h1;
  assign regs_368_clock = clock;
  assign regs_368_reset = reset;
  assign regs_369_io_in = 64'h0;
  assign regs_369_io_init = 64'h0;
  assign regs_369_io_enable = 1'h1;
  assign regs_369_clock = clock;
  assign regs_369_reset = reset;
  assign regs_370_io_in = 64'h0;
  assign regs_370_io_init = 64'h0;
  assign regs_370_io_enable = 1'h1;
  assign regs_370_clock = clock;
  assign regs_370_reset = reset;
  assign regs_371_io_in = 64'h0;
  assign regs_371_io_init = 64'h0;
  assign regs_371_io_enable = 1'h1;
  assign regs_371_clock = clock;
  assign regs_371_reset = reset;
  assign regs_372_io_in = 64'h0;
  assign regs_372_io_init = 64'h0;
  assign regs_372_io_enable = 1'h1;
  assign regs_372_clock = clock;
  assign regs_372_reset = reset;
  assign regs_373_io_in = 64'h0;
  assign regs_373_io_init = 64'h0;
  assign regs_373_io_enable = 1'h1;
  assign regs_373_clock = clock;
  assign regs_373_reset = reset;
  assign regs_374_io_in = 64'h0;
  assign regs_374_io_init = 64'h0;
  assign regs_374_io_enable = 1'h1;
  assign regs_374_clock = clock;
  assign regs_374_reset = reset;
  assign regs_375_io_in = 64'h0;
  assign regs_375_io_init = 64'h0;
  assign regs_375_io_enable = 1'h1;
  assign regs_375_clock = clock;
  assign regs_375_reset = reset;
  assign regs_376_io_in = 64'h0;
  assign regs_376_io_init = 64'h0;
  assign regs_376_io_enable = 1'h1;
  assign regs_376_clock = clock;
  assign regs_376_reset = reset;
  assign regs_377_io_in = 64'h0;
  assign regs_377_io_init = 64'h0;
  assign regs_377_io_enable = 1'h1;
  assign regs_377_clock = clock;
  assign regs_377_reset = reset;
  assign regs_378_io_in = 64'h0;
  assign regs_378_io_init = 64'h0;
  assign regs_378_io_enable = 1'h1;
  assign regs_378_clock = clock;
  assign regs_378_reset = reset;
  assign regs_379_io_in = 64'h0;
  assign regs_379_io_init = 64'h0;
  assign regs_379_io_enable = 1'h1;
  assign regs_379_clock = clock;
  assign regs_379_reset = reset;
  assign regs_380_io_in = 64'h0;
  assign regs_380_io_init = 64'h0;
  assign regs_380_io_enable = 1'h1;
  assign regs_380_clock = clock;
  assign regs_380_reset = reset;
  assign regs_381_io_in = 64'h0;
  assign regs_381_io_init = 64'h0;
  assign regs_381_io_enable = 1'h1;
  assign regs_381_clock = clock;
  assign regs_381_reset = reset;
  assign regs_382_io_in = 64'h0;
  assign regs_382_io_init = 64'h0;
  assign regs_382_io_enable = 1'h1;
  assign regs_382_clock = clock;
  assign regs_382_reset = reset;
  assign regs_383_io_in = 64'h0;
  assign regs_383_io_init = 64'h0;
  assign regs_383_io_enable = 1'h1;
  assign regs_383_clock = clock;
  assign regs_383_reset = reset;
  assign regs_384_io_in = 64'h0;
  assign regs_384_io_init = 64'h0;
  assign regs_384_io_enable = 1'h1;
  assign regs_384_clock = clock;
  assign regs_384_reset = reset;
  assign regs_385_io_in = 64'h0;
  assign regs_385_io_init = 64'h0;
  assign regs_385_io_enable = 1'h1;
  assign regs_385_clock = clock;
  assign regs_385_reset = reset;
  assign regs_386_io_in = 64'h0;
  assign regs_386_io_init = 64'h0;
  assign regs_386_io_enable = 1'h1;
  assign regs_386_clock = clock;
  assign regs_386_reset = reset;
  assign regs_387_io_in = 64'h0;
  assign regs_387_io_init = 64'h0;
  assign regs_387_io_enable = 1'h1;
  assign regs_387_clock = clock;
  assign regs_387_reset = reset;
  assign regs_388_io_in = 64'h0;
  assign regs_388_io_init = 64'h0;
  assign regs_388_io_enable = 1'h1;
  assign regs_388_clock = clock;
  assign regs_388_reset = reset;
  assign regs_389_io_in = 64'h0;
  assign regs_389_io_init = 64'h0;
  assign regs_389_io_enable = 1'h1;
  assign regs_389_clock = clock;
  assign regs_389_reset = reset;
  assign regs_390_io_in = 64'h0;
  assign regs_390_io_init = 64'h0;
  assign regs_390_io_enable = 1'h1;
  assign regs_390_clock = clock;
  assign regs_390_reset = reset;
  assign regs_391_io_in = 64'h0;
  assign regs_391_io_init = 64'h0;
  assign regs_391_io_enable = 1'h1;
  assign regs_391_clock = clock;
  assign regs_391_reset = reset;
  assign regs_392_io_in = 64'h0;
  assign regs_392_io_init = 64'h0;
  assign regs_392_io_enable = 1'h1;
  assign regs_392_clock = clock;
  assign regs_392_reset = reset;
  assign regs_393_io_in = 64'h0;
  assign regs_393_io_init = 64'h0;
  assign regs_393_io_enable = 1'h1;
  assign regs_393_clock = clock;
  assign regs_393_reset = reset;
  assign regs_394_io_in = 64'h0;
  assign regs_394_io_init = 64'h0;
  assign regs_394_io_enable = 1'h1;
  assign regs_394_clock = clock;
  assign regs_394_reset = reset;
  assign regs_395_io_in = 64'h0;
  assign regs_395_io_init = 64'h0;
  assign regs_395_io_enable = 1'h1;
  assign regs_395_clock = clock;
  assign regs_395_reset = reset;
  assign regs_396_io_in = 64'h0;
  assign regs_396_io_init = 64'h0;
  assign regs_396_io_enable = 1'h1;
  assign regs_396_clock = clock;
  assign regs_396_reset = reset;
  assign regs_397_io_in = 64'h0;
  assign regs_397_io_init = 64'h0;
  assign regs_397_io_enable = 1'h1;
  assign regs_397_clock = clock;
  assign regs_397_reset = reset;
  assign regs_398_io_in = 64'h0;
  assign regs_398_io_init = 64'h0;
  assign regs_398_io_enable = 1'h1;
  assign regs_398_clock = clock;
  assign regs_398_reset = reset;
  assign regs_399_io_in = 64'h0;
  assign regs_399_io_init = 64'h0;
  assign regs_399_io_enable = 1'h1;
  assign regs_399_clock = clock;
  assign regs_399_reset = reset;
  assign regs_400_io_in = 64'h0;
  assign regs_400_io_init = 64'h0;
  assign regs_400_io_enable = 1'h1;
  assign regs_400_clock = clock;
  assign regs_400_reset = reset;
  assign regs_401_io_in = 64'h0;
  assign regs_401_io_init = 64'h0;
  assign regs_401_io_enable = 1'h1;
  assign regs_401_clock = clock;
  assign regs_401_reset = reset;
  assign regs_402_io_in = 64'h0;
  assign regs_402_io_init = 64'h0;
  assign regs_402_io_enable = 1'h1;
  assign regs_402_clock = clock;
  assign regs_402_reset = reset;
  assign regs_403_io_in = 64'h0;
  assign regs_403_io_init = 64'h0;
  assign regs_403_io_enable = 1'h1;
  assign regs_403_clock = clock;
  assign regs_403_reset = reset;
  assign regs_404_io_in = 64'h0;
  assign regs_404_io_init = 64'h0;
  assign regs_404_io_enable = 1'h1;
  assign regs_404_clock = clock;
  assign regs_404_reset = reset;
  assign regs_405_io_in = 64'h0;
  assign regs_405_io_init = 64'h0;
  assign regs_405_io_enable = 1'h1;
  assign regs_405_clock = clock;
  assign regs_405_reset = reset;
  assign regs_406_io_in = 64'h0;
  assign regs_406_io_init = 64'h0;
  assign regs_406_io_enable = 1'h1;
  assign regs_406_clock = clock;
  assign regs_406_reset = reset;
  assign regs_407_io_in = 64'h0;
  assign regs_407_io_init = 64'h0;
  assign regs_407_io_enable = 1'h1;
  assign regs_407_clock = clock;
  assign regs_407_reset = reset;
  assign regs_408_io_in = 64'h0;
  assign regs_408_io_init = 64'h0;
  assign regs_408_io_enable = 1'h1;
  assign regs_408_clock = clock;
  assign regs_408_reset = reset;
  assign regs_409_io_in = 64'h0;
  assign regs_409_io_init = 64'h0;
  assign regs_409_io_enable = 1'h1;
  assign regs_409_clock = clock;
  assign regs_409_reset = reset;
  assign regs_410_io_in = 64'h0;
  assign regs_410_io_init = 64'h0;
  assign regs_410_io_enable = 1'h1;
  assign regs_410_clock = clock;
  assign regs_410_reset = reset;
  assign regs_411_io_in = 64'h0;
  assign regs_411_io_init = 64'h0;
  assign regs_411_io_enable = 1'h1;
  assign regs_411_clock = clock;
  assign regs_411_reset = reset;
  assign regs_412_io_in = 64'h0;
  assign regs_412_io_init = 64'h0;
  assign regs_412_io_enable = 1'h1;
  assign regs_412_clock = clock;
  assign regs_412_reset = reset;
  assign regs_413_io_in = 64'h0;
  assign regs_413_io_init = 64'h0;
  assign regs_413_io_enable = 1'h1;
  assign regs_413_clock = clock;
  assign regs_413_reset = reset;
  assign regs_414_io_in = 64'h0;
  assign regs_414_io_init = 64'h0;
  assign regs_414_io_enable = 1'h1;
  assign regs_414_clock = clock;
  assign regs_414_reset = reset;
  assign regs_415_io_in = 64'h0;
  assign regs_415_io_init = 64'h0;
  assign regs_415_io_enable = 1'h1;
  assign regs_415_clock = clock;
  assign regs_415_reset = reset;
  assign regs_416_io_in = 64'h0;
  assign regs_416_io_init = 64'h0;
  assign regs_416_io_enable = 1'h1;
  assign regs_416_clock = clock;
  assign regs_416_reset = reset;
  assign regs_417_io_in = 64'h0;
  assign regs_417_io_init = 64'h0;
  assign regs_417_io_enable = 1'h1;
  assign regs_417_clock = clock;
  assign regs_417_reset = reset;
  assign regs_418_io_in = 64'h0;
  assign regs_418_io_init = 64'h0;
  assign regs_418_io_enable = 1'h1;
  assign regs_418_clock = clock;
  assign regs_418_reset = reset;
  assign regs_419_io_in = 64'h0;
  assign regs_419_io_init = 64'h0;
  assign regs_419_io_enable = 1'h1;
  assign regs_419_clock = clock;
  assign regs_419_reset = reset;
  assign regs_420_io_in = 64'h0;
  assign regs_420_io_init = 64'h0;
  assign regs_420_io_enable = 1'h1;
  assign regs_420_clock = clock;
  assign regs_420_reset = reset;
  assign regs_421_io_in = 64'h0;
  assign regs_421_io_init = 64'h0;
  assign regs_421_io_enable = 1'h1;
  assign regs_421_clock = clock;
  assign regs_421_reset = reset;
  assign regs_422_io_in = 64'h0;
  assign regs_422_io_init = 64'h0;
  assign regs_422_io_enable = 1'h1;
  assign regs_422_clock = clock;
  assign regs_422_reset = reset;
  assign regs_423_io_in = 64'h0;
  assign regs_423_io_init = 64'h0;
  assign regs_423_io_enable = 1'h1;
  assign regs_423_clock = clock;
  assign regs_423_reset = reset;
  assign regs_424_io_in = 64'h0;
  assign regs_424_io_init = 64'h0;
  assign regs_424_io_enable = 1'h1;
  assign regs_424_clock = clock;
  assign regs_424_reset = reset;
  assign regs_425_io_in = 64'h0;
  assign regs_425_io_init = 64'h0;
  assign regs_425_io_enable = 1'h1;
  assign regs_425_clock = clock;
  assign regs_425_reset = reset;
  assign regs_426_io_in = 64'h0;
  assign regs_426_io_init = 64'h0;
  assign regs_426_io_enable = 1'h1;
  assign regs_426_clock = clock;
  assign regs_426_reset = reset;
  assign regs_427_io_in = 64'h0;
  assign regs_427_io_init = 64'h0;
  assign regs_427_io_enable = 1'h1;
  assign regs_427_clock = clock;
  assign regs_427_reset = reset;
  assign regs_428_io_in = 64'h0;
  assign regs_428_io_init = 64'h0;
  assign regs_428_io_enable = 1'h1;
  assign regs_428_clock = clock;
  assign regs_428_reset = reset;
  assign regs_429_io_in = 64'h0;
  assign regs_429_io_init = 64'h0;
  assign regs_429_io_enable = 1'h1;
  assign regs_429_clock = clock;
  assign regs_429_reset = reset;
  assign regs_430_io_in = 64'h0;
  assign regs_430_io_init = 64'h0;
  assign regs_430_io_enable = 1'h1;
  assign regs_430_clock = clock;
  assign regs_430_reset = reset;
  assign regs_431_io_in = 64'h0;
  assign regs_431_io_init = 64'h0;
  assign regs_431_io_enable = 1'h1;
  assign regs_431_clock = clock;
  assign regs_431_reset = reset;
  assign regs_432_io_in = 64'h0;
  assign regs_432_io_init = 64'h0;
  assign regs_432_io_enable = 1'h1;
  assign regs_432_clock = clock;
  assign regs_432_reset = reset;
  assign regs_433_io_in = 64'h0;
  assign regs_433_io_init = 64'h0;
  assign regs_433_io_enable = 1'h1;
  assign regs_433_clock = clock;
  assign regs_433_reset = reset;
  assign regs_434_io_in = 64'h0;
  assign regs_434_io_init = 64'h0;
  assign regs_434_io_enable = 1'h1;
  assign regs_434_clock = clock;
  assign regs_434_reset = reset;
  assign regs_435_io_in = 64'h0;
  assign regs_435_io_init = 64'h0;
  assign regs_435_io_enable = 1'h1;
  assign regs_435_clock = clock;
  assign regs_435_reset = reset;
  assign regs_436_io_in = 64'h0;
  assign regs_436_io_init = 64'h0;
  assign regs_436_io_enable = 1'h1;
  assign regs_436_clock = clock;
  assign regs_436_reset = reset;
  assign regs_437_io_in = 64'h0;
  assign regs_437_io_init = 64'h0;
  assign regs_437_io_enable = 1'h1;
  assign regs_437_clock = clock;
  assign regs_437_reset = reset;
  assign regs_438_io_in = 64'h0;
  assign regs_438_io_init = 64'h0;
  assign regs_438_io_enable = 1'h1;
  assign regs_438_clock = clock;
  assign regs_438_reset = reset;
  assign regs_439_io_in = 64'h0;
  assign regs_439_io_init = 64'h0;
  assign regs_439_io_enable = 1'h1;
  assign regs_439_clock = clock;
  assign regs_439_reset = reset;
  assign regs_440_io_in = 64'h0;
  assign regs_440_io_init = 64'h0;
  assign regs_440_io_enable = 1'h1;
  assign regs_440_clock = clock;
  assign regs_440_reset = reset;
  assign regs_441_io_in = 64'h0;
  assign regs_441_io_init = 64'h0;
  assign regs_441_io_enable = 1'h1;
  assign regs_441_clock = clock;
  assign regs_441_reset = reset;
  assign regs_442_io_in = 64'h0;
  assign regs_442_io_init = 64'h0;
  assign regs_442_io_enable = 1'h1;
  assign regs_442_clock = clock;
  assign regs_442_reset = reset;
  assign regs_443_io_in = 64'h0;
  assign regs_443_io_init = 64'h0;
  assign regs_443_io_enable = 1'h1;
  assign regs_443_clock = clock;
  assign regs_443_reset = reset;
  assign regs_444_io_in = 64'h0;
  assign regs_444_io_init = 64'h0;
  assign regs_444_io_enable = 1'h1;
  assign regs_444_clock = clock;
  assign regs_444_reset = reset;
  assign regs_445_io_in = 64'h0;
  assign regs_445_io_init = 64'h0;
  assign regs_445_io_enable = 1'h1;
  assign regs_445_clock = clock;
  assign regs_445_reset = reset;
  assign regs_446_io_in = 64'h0;
  assign regs_446_io_init = 64'h0;
  assign regs_446_io_enable = 1'h1;
  assign regs_446_clock = clock;
  assign regs_446_reset = reset;
  assign regs_447_io_in = 64'h0;
  assign regs_447_io_init = 64'h0;
  assign regs_447_io_enable = 1'h1;
  assign regs_447_clock = clock;
  assign regs_447_reset = reset;
  assign regs_448_io_in = 64'h0;
  assign regs_448_io_init = 64'h0;
  assign regs_448_io_enable = 1'h1;
  assign regs_448_clock = clock;
  assign regs_448_reset = reset;
  assign regs_449_io_in = 64'h0;
  assign regs_449_io_init = 64'h0;
  assign regs_449_io_enable = 1'h1;
  assign regs_449_clock = clock;
  assign regs_449_reset = reset;
  assign regs_450_io_in = 64'h0;
  assign regs_450_io_init = 64'h0;
  assign regs_450_io_enable = 1'h1;
  assign regs_450_clock = clock;
  assign regs_450_reset = reset;
  assign regs_451_io_in = 64'h0;
  assign regs_451_io_init = 64'h0;
  assign regs_451_io_enable = 1'h1;
  assign regs_451_clock = clock;
  assign regs_451_reset = reset;
  assign regs_452_io_in = 64'h0;
  assign regs_452_io_init = 64'h0;
  assign regs_452_io_enable = 1'h1;
  assign regs_452_clock = clock;
  assign regs_452_reset = reset;
  assign regs_453_io_in = 64'h0;
  assign regs_453_io_init = 64'h0;
  assign regs_453_io_enable = 1'h1;
  assign regs_453_clock = clock;
  assign regs_453_reset = reset;
  assign regs_454_io_in = 64'h0;
  assign regs_454_io_init = 64'h0;
  assign regs_454_io_enable = 1'h1;
  assign regs_454_clock = clock;
  assign regs_454_reset = reset;
  assign regs_455_io_in = 64'h0;
  assign regs_455_io_init = 64'h0;
  assign regs_455_io_enable = 1'h1;
  assign regs_455_clock = clock;
  assign regs_455_reset = reset;
  assign regs_456_io_in = 64'h0;
  assign regs_456_io_init = 64'h0;
  assign regs_456_io_enable = 1'h1;
  assign regs_456_clock = clock;
  assign regs_456_reset = reset;
  assign regs_457_io_in = 64'h0;
  assign regs_457_io_init = 64'h0;
  assign regs_457_io_enable = 1'h1;
  assign regs_457_clock = clock;
  assign regs_457_reset = reset;
  assign regs_458_io_in = 64'h0;
  assign regs_458_io_init = 64'h0;
  assign regs_458_io_enable = 1'h1;
  assign regs_458_clock = clock;
  assign regs_458_reset = reset;
  assign regs_459_io_in = 64'h0;
  assign regs_459_io_init = 64'h0;
  assign regs_459_io_enable = 1'h1;
  assign regs_459_clock = clock;
  assign regs_459_reset = reset;
  assign regs_460_io_in = 64'h0;
  assign regs_460_io_init = 64'h0;
  assign regs_460_io_enable = 1'h1;
  assign regs_460_clock = clock;
  assign regs_460_reset = reset;
  assign regs_461_io_in = 64'h0;
  assign regs_461_io_init = 64'h0;
  assign regs_461_io_enable = 1'h1;
  assign regs_461_clock = clock;
  assign regs_461_reset = reset;
  assign regs_462_io_in = 64'h0;
  assign regs_462_io_init = 64'h0;
  assign regs_462_io_enable = 1'h1;
  assign regs_462_clock = clock;
  assign regs_462_reset = reset;
  assign regs_463_io_in = 64'h0;
  assign regs_463_io_init = 64'h0;
  assign regs_463_io_enable = 1'h1;
  assign regs_463_clock = clock;
  assign regs_463_reset = reset;
  assign regs_464_io_in = 64'h0;
  assign regs_464_io_init = 64'h0;
  assign regs_464_io_enable = 1'h1;
  assign regs_464_clock = clock;
  assign regs_464_reset = reset;
  assign regs_465_io_in = 64'h0;
  assign regs_465_io_init = 64'h0;
  assign regs_465_io_enable = 1'h1;
  assign regs_465_clock = clock;
  assign regs_465_reset = reset;
  assign regs_466_io_in = 64'h0;
  assign regs_466_io_init = 64'h0;
  assign regs_466_io_enable = 1'h1;
  assign regs_466_clock = clock;
  assign regs_466_reset = reset;
  assign regs_467_io_in = 64'h0;
  assign regs_467_io_init = 64'h0;
  assign regs_467_io_enable = 1'h1;
  assign regs_467_clock = clock;
  assign regs_467_reset = reset;
  assign regs_468_io_in = 64'h0;
  assign regs_468_io_init = 64'h0;
  assign regs_468_io_enable = 1'h1;
  assign regs_468_clock = clock;
  assign regs_468_reset = reset;
  assign regs_469_io_in = 64'h0;
  assign regs_469_io_init = 64'h0;
  assign regs_469_io_enable = 1'h1;
  assign regs_469_clock = clock;
  assign regs_469_reset = reset;
  assign regs_470_io_in = 64'h0;
  assign regs_470_io_init = 64'h0;
  assign regs_470_io_enable = 1'h1;
  assign regs_470_clock = clock;
  assign regs_470_reset = reset;
  assign regs_471_io_in = 64'h0;
  assign regs_471_io_init = 64'h0;
  assign regs_471_io_enable = 1'h1;
  assign regs_471_clock = clock;
  assign regs_471_reset = reset;
  assign regs_472_io_in = 64'h0;
  assign regs_472_io_init = 64'h0;
  assign regs_472_io_enable = 1'h1;
  assign regs_472_clock = clock;
  assign regs_472_reset = reset;
  assign regs_473_io_in = 64'h0;
  assign regs_473_io_init = 64'h0;
  assign regs_473_io_enable = 1'h1;
  assign regs_473_clock = clock;
  assign regs_473_reset = reset;
  assign regs_474_io_in = 64'h0;
  assign regs_474_io_init = 64'h0;
  assign regs_474_io_enable = 1'h1;
  assign regs_474_clock = clock;
  assign regs_474_reset = reset;
  assign regs_475_io_in = 64'h0;
  assign regs_475_io_init = 64'h0;
  assign regs_475_io_enable = 1'h1;
  assign regs_475_clock = clock;
  assign regs_475_reset = reset;
  assign regs_476_io_in = 64'h0;
  assign regs_476_io_init = 64'h0;
  assign regs_476_io_enable = 1'h1;
  assign regs_476_clock = clock;
  assign regs_476_reset = reset;
  assign regs_477_io_in = 64'h0;
  assign regs_477_io_init = 64'h0;
  assign regs_477_io_enable = 1'h1;
  assign regs_477_clock = clock;
  assign regs_477_reset = reset;
  assign regs_478_io_in = 64'h0;
  assign regs_478_io_init = 64'h0;
  assign regs_478_io_enable = 1'h1;
  assign regs_478_clock = clock;
  assign regs_478_reset = reset;
  assign regs_479_io_in = 64'h0;
  assign regs_479_io_init = 64'h0;
  assign regs_479_io_enable = 1'h1;
  assign regs_479_clock = clock;
  assign regs_479_reset = reset;
  assign regs_480_io_in = 64'h0;
  assign regs_480_io_init = 64'h0;
  assign regs_480_io_enable = 1'h1;
  assign regs_480_clock = clock;
  assign regs_480_reset = reset;
  assign regs_481_io_in = 64'h0;
  assign regs_481_io_init = 64'h0;
  assign regs_481_io_enable = 1'h1;
  assign regs_481_clock = clock;
  assign regs_481_reset = reset;
  assign regs_482_io_in = 64'h0;
  assign regs_482_io_init = 64'h0;
  assign regs_482_io_enable = 1'h1;
  assign regs_482_clock = clock;
  assign regs_482_reset = reset;
  assign regs_483_io_in = 64'h0;
  assign regs_483_io_init = 64'h0;
  assign regs_483_io_enable = 1'h1;
  assign regs_483_clock = clock;
  assign regs_483_reset = reset;
  assign regs_484_io_in = 64'h0;
  assign regs_484_io_init = 64'h0;
  assign regs_484_io_enable = 1'h1;
  assign regs_484_clock = clock;
  assign regs_484_reset = reset;
  assign regs_485_io_in = 64'h0;
  assign regs_485_io_init = 64'h0;
  assign regs_485_io_enable = 1'h1;
  assign regs_485_clock = clock;
  assign regs_485_reset = reset;
  assign regs_486_io_in = 64'h0;
  assign regs_486_io_init = 64'h0;
  assign regs_486_io_enable = 1'h1;
  assign regs_486_clock = clock;
  assign regs_486_reset = reset;
  assign regs_487_io_in = 64'h0;
  assign regs_487_io_init = 64'h0;
  assign regs_487_io_enable = 1'h1;
  assign regs_487_clock = clock;
  assign regs_487_reset = reset;
  assign regs_488_io_in = 64'h0;
  assign regs_488_io_init = 64'h0;
  assign regs_488_io_enable = 1'h1;
  assign regs_488_clock = clock;
  assign regs_488_reset = reset;
  assign regs_489_io_in = 64'h0;
  assign regs_489_io_init = 64'h0;
  assign regs_489_io_enable = 1'h1;
  assign regs_489_clock = clock;
  assign regs_489_reset = reset;
  assign regs_490_io_in = 64'h0;
  assign regs_490_io_init = 64'h0;
  assign regs_490_io_enable = 1'h1;
  assign regs_490_clock = clock;
  assign regs_490_reset = reset;
  assign regs_491_io_in = 64'h0;
  assign regs_491_io_init = 64'h0;
  assign regs_491_io_enable = 1'h1;
  assign regs_491_clock = clock;
  assign regs_491_reset = reset;
  assign regs_492_io_in = 64'h0;
  assign regs_492_io_init = 64'h0;
  assign regs_492_io_enable = 1'h1;
  assign regs_492_clock = clock;
  assign regs_492_reset = reset;
  assign regs_493_io_in = 64'h0;
  assign regs_493_io_init = 64'h0;
  assign regs_493_io_enable = 1'h1;
  assign regs_493_clock = clock;
  assign regs_493_reset = reset;
  assign regs_494_io_in = 64'h0;
  assign regs_494_io_init = 64'h0;
  assign regs_494_io_enable = 1'h1;
  assign regs_494_clock = clock;
  assign regs_494_reset = reset;
  assign regs_495_io_in = 64'h0;
  assign regs_495_io_init = 64'h0;
  assign regs_495_io_enable = 1'h1;
  assign regs_495_clock = clock;
  assign regs_495_reset = reset;
  assign regs_496_io_in = 64'h0;
  assign regs_496_io_init = 64'h0;
  assign regs_496_io_enable = 1'h1;
  assign regs_496_clock = clock;
  assign regs_496_reset = reset;
  assign regs_497_io_in = 64'h0;
  assign regs_497_io_init = 64'h0;
  assign regs_497_io_enable = 1'h1;
  assign regs_497_clock = clock;
  assign regs_497_reset = reset;
  assign regs_498_io_in = 64'h0;
  assign regs_498_io_init = 64'h0;
  assign regs_498_io_enable = 1'h1;
  assign regs_498_clock = clock;
  assign regs_498_reset = reset;
  assign regs_499_io_in = 64'h0;
  assign regs_499_io_init = 64'h0;
  assign regs_499_io_enable = 1'h1;
  assign regs_499_clock = clock;
  assign regs_499_reset = reset;
  assign regs_500_io_in = 64'h0;
  assign regs_500_io_init = 64'h0;
  assign regs_500_io_enable = 1'h1;
  assign regs_500_clock = clock;
  assign regs_500_reset = reset;
  assign regs_501_io_in = 64'h0;
  assign regs_501_io_init = 64'h0;
  assign regs_501_io_enable = 1'h1;
  assign regs_501_clock = clock;
  assign regs_501_reset = reset;
  assign regs_502_io_in = 64'h0;
  assign regs_502_io_init = 64'h0;
  assign regs_502_io_enable = 1'h1;
  assign regs_502_clock = clock;
  assign regs_502_reset = reset;
  assign regs_503_io_in = 64'h0;
  assign regs_503_io_init = 64'h0;
  assign regs_503_io_enable = 1'h1;
  assign regs_503_clock = clock;
  assign regs_503_reset = reset;
  assign regs_504_io_in = 64'h0;
  assign regs_504_io_init = 64'h0;
  assign regs_504_io_enable = 1'h1;
  assign regs_504_clock = clock;
  assign regs_504_reset = reset;
  assign rport_io_ins_0 = regOuts_0;
  assign rport_io_ins_1 = regOuts_1;
  assign rport_io_ins_2 = regOuts_2;
  assign rport_io_ins_3 = regOuts_3;
  assign rport_io_ins_4 = regOuts_4;
  assign rport_io_ins_5 = regOuts_5;
  assign rport_io_ins_6 = regOuts_6;
  assign rport_io_ins_7 = regOuts_7;
  assign rport_io_ins_8 = regOuts_8;
  assign rport_io_ins_9 = regOuts_9;
  assign rport_io_ins_10 = regOuts_10;
  assign rport_io_ins_11 = regOuts_11;
  assign rport_io_ins_12 = regOuts_12;
  assign rport_io_ins_13 = regOuts_13;
  assign rport_io_ins_14 = regOuts_14;
  assign rport_io_ins_15 = regOuts_15;
  assign rport_io_ins_16 = regOuts_16;
  assign rport_io_ins_17 = regOuts_17;
  assign rport_io_ins_18 = regOuts_18;
  assign rport_io_ins_19 = regOuts_19;
  assign rport_io_ins_20 = regOuts_20;
  assign rport_io_ins_21 = regOuts_21;
  assign rport_io_ins_22 = regOuts_22;
  assign rport_io_ins_23 = regOuts_23;
  assign rport_io_ins_24 = regOuts_24;
  assign rport_io_ins_25 = regOuts_25;
  assign rport_io_ins_26 = regOuts_26;
  assign rport_io_ins_27 = regOuts_27;
  assign rport_io_ins_28 = regOuts_28;
  assign rport_io_ins_29 = regOuts_29;
  assign rport_io_ins_30 = regOuts_30;
  assign rport_io_ins_31 = regOuts_31;
  assign rport_io_ins_32 = regOuts_32;
  assign rport_io_ins_33 = regOuts_33;
  assign rport_io_ins_34 = regOuts_34;
  assign rport_io_ins_35 = regOuts_35;
  assign rport_io_ins_36 = regOuts_36;
  assign rport_io_ins_37 = regOuts_37;
  assign rport_io_ins_38 = regOuts_38;
  assign rport_io_ins_39 = regOuts_39;
  assign rport_io_ins_40 = regOuts_40;
  assign rport_io_ins_41 = regOuts_41;
  assign rport_io_ins_42 = regOuts_42;
  assign rport_io_ins_43 = regOuts_43;
  assign rport_io_ins_44 = regOuts_44;
  assign rport_io_ins_45 = regOuts_45;
  assign rport_io_ins_46 = regOuts_46;
  assign rport_io_ins_47 = regOuts_47;
  assign rport_io_ins_48 = regOuts_48;
  assign rport_io_ins_49 = regOuts_49;
  assign rport_io_ins_50 = regOuts_50;
  assign rport_io_ins_51 = regOuts_51;
  assign rport_io_ins_52 = regOuts_52;
  assign rport_io_ins_53 = regOuts_53;
  assign rport_io_ins_54 = regOuts_54;
  assign rport_io_ins_55 = regOuts_55;
  assign rport_io_ins_56 = regOuts_56;
  assign rport_io_ins_57 = regOuts_57;
  assign rport_io_ins_58 = regOuts_58;
  assign rport_io_ins_59 = regOuts_59;
  assign rport_io_ins_60 = regOuts_60;
  assign rport_io_ins_61 = regOuts_61;
  assign rport_io_ins_62 = regOuts_62;
  assign rport_io_ins_63 = regOuts_63;
  assign rport_io_ins_64 = regOuts_64;
  assign rport_io_ins_65 = regOuts_65;
  assign rport_io_ins_66 = regOuts_66;
  assign rport_io_ins_67 = regOuts_67;
  assign rport_io_ins_68 = regOuts_68;
  assign rport_io_ins_69 = regOuts_69;
  assign rport_io_ins_70 = regOuts_70;
  assign rport_io_ins_71 = regOuts_71;
  assign rport_io_ins_72 = regOuts_72;
  assign rport_io_ins_73 = regOuts_73;
  assign rport_io_ins_74 = regOuts_74;
  assign rport_io_ins_75 = regOuts_75;
  assign rport_io_ins_76 = regOuts_76;
  assign rport_io_ins_77 = regOuts_77;
  assign rport_io_ins_78 = regOuts_78;
  assign rport_io_ins_79 = regOuts_79;
  assign rport_io_ins_80 = regOuts_80;
  assign rport_io_ins_81 = regOuts_81;
  assign rport_io_ins_82 = regOuts_82;
  assign rport_io_ins_83 = regOuts_83;
  assign rport_io_ins_84 = regOuts_84;
  assign rport_io_ins_85 = regOuts_85;
  assign rport_io_ins_86 = regOuts_86;
  assign rport_io_ins_87 = regOuts_87;
  assign rport_io_ins_88 = regOuts_88;
  assign rport_io_ins_89 = regOuts_89;
  assign rport_io_ins_90 = regOuts_90;
  assign rport_io_ins_91 = regOuts_91;
  assign rport_io_ins_92 = regOuts_92;
  assign rport_io_ins_93 = regOuts_93;
  assign rport_io_ins_94 = regOuts_94;
  assign rport_io_ins_95 = regOuts_95;
  assign rport_io_ins_96 = regOuts_96;
  assign rport_io_ins_97 = regOuts_97;
  assign rport_io_ins_98 = regOuts_98;
  assign rport_io_ins_99 = regOuts_99;
  assign rport_io_ins_100 = regOuts_100;
  assign rport_io_ins_101 = regOuts_101;
  assign rport_io_ins_102 = regOuts_102;
  assign rport_io_ins_103 = regOuts_103;
  assign rport_io_ins_104 = regOuts_104;
  assign rport_io_ins_105 = regOuts_105;
  assign rport_io_ins_106 = regOuts_106;
  assign rport_io_ins_107 = regOuts_107;
  assign rport_io_ins_108 = regOuts_108;
  assign rport_io_ins_109 = regOuts_109;
  assign rport_io_ins_110 = regOuts_110;
  assign rport_io_ins_111 = regOuts_111;
  assign rport_io_ins_112 = regOuts_112;
  assign rport_io_ins_113 = regOuts_113;
  assign rport_io_ins_114 = regOuts_114;
  assign rport_io_ins_115 = regOuts_115;
  assign rport_io_ins_116 = regOuts_116;
  assign rport_io_ins_117 = regOuts_117;
  assign rport_io_ins_118 = regOuts_118;
  assign rport_io_ins_119 = regOuts_119;
  assign rport_io_ins_120 = regOuts_120;
  assign rport_io_ins_121 = regOuts_121;
  assign rport_io_ins_122 = regOuts_122;
  assign rport_io_ins_123 = regOuts_123;
  assign rport_io_ins_124 = regOuts_124;
  assign rport_io_ins_125 = regOuts_125;
  assign rport_io_ins_126 = regOuts_126;
  assign rport_io_ins_127 = regOuts_127;
  assign rport_io_ins_128 = regOuts_128;
  assign rport_io_ins_129 = regOuts_129;
  assign rport_io_ins_130 = regOuts_130;
  assign rport_io_ins_131 = regOuts_131;
  assign rport_io_ins_132 = regOuts_132;
  assign rport_io_ins_133 = regOuts_133;
  assign rport_io_ins_134 = regOuts_134;
  assign rport_io_ins_135 = regOuts_135;
  assign rport_io_ins_136 = regOuts_136;
  assign rport_io_ins_137 = regOuts_137;
  assign rport_io_ins_138 = regOuts_138;
  assign rport_io_ins_139 = regOuts_139;
  assign rport_io_ins_140 = regOuts_140;
  assign rport_io_ins_141 = regOuts_141;
  assign rport_io_ins_142 = regOuts_142;
  assign rport_io_ins_143 = regOuts_143;
  assign rport_io_ins_144 = regOuts_144;
  assign rport_io_ins_145 = regOuts_145;
  assign rport_io_ins_146 = regOuts_146;
  assign rport_io_ins_147 = regOuts_147;
  assign rport_io_ins_148 = regOuts_148;
  assign rport_io_ins_149 = regOuts_149;
  assign rport_io_ins_150 = regOuts_150;
  assign rport_io_ins_151 = regOuts_151;
  assign rport_io_ins_152 = regOuts_152;
  assign rport_io_ins_153 = regOuts_153;
  assign rport_io_ins_154 = regOuts_154;
  assign rport_io_ins_155 = regOuts_155;
  assign rport_io_ins_156 = regOuts_156;
  assign rport_io_ins_157 = regOuts_157;
  assign rport_io_ins_158 = regOuts_158;
  assign rport_io_ins_159 = regOuts_159;
  assign rport_io_ins_160 = regOuts_160;
  assign rport_io_ins_161 = regOuts_161;
  assign rport_io_ins_162 = regOuts_162;
  assign rport_io_ins_163 = regOuts_163;
  assign rport_io_ins_164 = regOuts_164;
  assign rport_io_ins_165 = regOuts_165;
  assign rport_io_ins_166 = regOuts_166;
  assign rport_io_ins_167 = regOuts_167;
  assign rport_io_ins_168 = regOuts_168;
  assign rport_io_ins_169 = regOuts_169;
  assign rport_io_ins_170 = regOuts_170;
  assign rport_io_ins_171 = regOuts_171;
  assign rport_io_ins_172 = regOuts_172;
  assign rport_io_ins_173 = regOuts_173;
  assign rport_io_ins_174 = regOuts_174;
  assign rport_io_ins_175 = regOuts_175;
  assign rport_io_ins_176 = regOuts_176;
  assign rport_io_ins_177 = regOuts_177;
  assign rport_io_ins_178 = regOuts_178;
  assign rport_io_ins_179 = regOuts_179;
  assign rport_io_ins_180 = regOuts_180;
  assign rport_io_ins_181 = regOuts_181;
  assign rport_io_ins_182 = regOuts_182;
  assign rport_io_ins_183 = regOuts_183;
  assign rport_io_ins_184 = regOuts_184;
  assign rport_io_ins_185 = regOuts_185;
  assign rport_io_ins_186 = regOuts_186;
  assign rport_io_ins_187 = regOuts_187;
  assign rport_io_ins_188 = regOuts_188;
  assign rport_io_ins_189 = regOuts_189;
  assign rport_io_ins_190 = regOuts_190;
  assign rport_io_ins_191 = regOuts_191;
  assign rport_io_ins_192 = regOuts_192;
  assign rport_io_ins_193 = regOuts_193;
  assign rport_io_ins_194 = regOuts_194;
  assign rport_io_ins_195 = regOuts_195;
  assign rport_io_ins_196 = regOuts_196;
  assign rport_io_ins_197 = regOuts_197;
  assign rport_io_ins_198 = regOuts_198;
  assign rport_io_ins_199 = regOuts_199;
  assign rport_io_ins_200 = regOuts_200;
  assign rport_io_ins_201 = regOuts_201;
  assign rport_io_ins_202 = regOuts_202;
  assign rport_io_ins_203 = regOuts_203;
  assign rport_io_ins_204 = regOuts_204;
  assign rport_io_ins_205 = regOuts_205;
  assign rport_io_ins_206 = regOuts_206;
  assign rport_io_ins_207 = regOuts_207;
  assign rport_io_ins_208 = regOuts_208;
  assign rport_io_ins_209 = regOuts_209;
  assign rport_io_ins_210 = regOuts_210;
  assign rport_io_ins_211 = regOuts_211;
  assign rport_io_ins_212 = regOuts_212;
  assign rport_io_ins_213 = regOuts_213;
  assign rport_io_ins_214 = regOuts_214;
  assign rport_io_ins_215 = regOuts_215;
  assign rport_io_ins_216 = regOuts_216;
  assign rport_io_ins_217 = regOuts_217;
  assign rport_io_ins_218 = regOuts_218;
  assign rport_io_ins_219 = regOuts_219;
  assign rport_io_ins_220 = regOuts_220;
  assign rport_io_ins_221 = regOuts_221;
  assign rport_io_ins_222 = regOuts_222;
  assign rport_io_ins_223 = regOuts_223;
  assign rport_io_ins_224 = regOuts_224;
  assign rport_io_ins_225 = regOuts_225;
  assign rport_io_ins_226 = regOuts_226;
  assign rport_io_ins_227 = regOuts_227;
  assign rport_io_ins_228 = regOuts_228;
  assign rport_io_ins_229 = regOuts_229;
  assign rport_io_ins_230 = regOuts_230;
  assign rport_io_ins_231 = regOuts_231;
  assign rport_io_ins_232 = regOuts_232;
  assign rport_io_ins_233 = regOuts_233;
  assign rport_io_ins_234 = regOuts_234;
  assign rport_io_ins_235 = regOuts_235;
  assign rport_io_ins_236 = regOuts_236;
  assign rport_io_ins_237 = regOuts_237;
  assign rport_io_ins_238 = regOuts_238;
  assign rport_io_ins_239 = regOuts_239;
  assign rport_io_ins_240 = regOuts_240;
  assign rport_io_ins_241 = regOuts_241;
  assign rport_io_ins_242 = regOuts_242;
  assign rport_io_ins_243 = regOuts_243;
  assign rport_io_ins_244 = regOuts_244;
  assign rport_io_ins_245 = regOuts_245;
  assign rport_io_ins_246 = regOuts_246;
  assign rport_io_ins_247 = regOuts_247;
  assign rport_io_ins_248 = regOuts_248;
  assign rport_io_ins_249 = regOuts_249;
  assign rport_io_ins_250 = regOuts_250;
  assign rport_io_ins_251 = regOuts_251;
  assign rport_io_ins_252 = regOuts_252;
  assign rport_io_ins_253 = regOuts_253;
  assign rport_io_ins_254 = regOuts_254;
  assign rport_io_ins_255 = regOuts_255;
  assign rport_io_ins_256 = regOuts_256;
  assign rport_io_ins_257 = regOuts_257;
  assign rport_io_ins_258 = regOuts_258;
  assign rport_io_ins_259 = regOuts_259;
  assign rport_io_ins_260 = regOuts_260;
  assign rport_io_ins_261 = regOuts_261;
  assign rport_io_ins_262 = regOuts_262;
  assign rport_io_ins_263 = regOuts_263;
  assign rport_io_ins_264 = regOuts_264;
  assign rport_io_ins_265 = regOuts_265;
  assign rport_io_ins_266 = regOuts_266;
  assign rport_io_ins_267 = regOuts_267;
  assign rport_io_ins_268 = regOuts_268;
  assign rport_io_ins_269 = regOuts_269;
  assign rport_io_ins_270 = regOuts_270;
  assign rport_io_ins_271 = regOuts_271;
  assign rport_io_ins_272 = regOuts_272;
  assign rport_io_ins_273 = regOuts_273;
  assign rport_io_ins_274 = regOuts_274;
  assign rport_io_ins_275 = regOuts_275;
  assign rport_io_ins_276 = regOuts_276;
  assign rport_io_ins_277 = regOuts_277;
  assign rport_io_ins_278 = regOuts_278;
  assign rport_io_ins_279 = regOuts_279;
  assign rport_io_ins_280 = regOuts_280;
  assign rport_io_ins_281 = regOuts_281;
  assign rport_io_ins_282 = regOuts_282;
  assign rport_io_ins_283 = regOuts_283;
  assign rport_io_ins_284 = regOuts_284;
  assign rport_io_ins_285 = regOuts_285;
  assign rport_io_ins_286 = regOuts_286;
  assign rport_io_ins_287 = regOuts_287;
  assign rport_io_ins_288 = regOuts_288;
  assign rport_io_ins_289 = regOuts_289;
  assign rport_io_ins_290 = regOuts_290;
  assign rport_io_ins_291 = regOuts_291;
  assign rport_io_ins_292 = regOuts_292;
  assign rport_io_ins_293 = regOuts_293;
  assign rport_io_ins_294 = regOuts_294;
  assign rport_io_ins_295 = regOuts_295;
  assign rport_io_ins_296 = regOuts_296;
  assign rport_io_ins_297 = regOuts_297;
  assign rport_io_ins_298 = regOuts_298;
  assign rport_io_ins_299 = regOuts_299;
  assign rport_io_ins_300 = regOuts_300;
  assign rport_io_ins_301 = regOuts_301;
  assign rport_io_ins_302 = regOuts_302;
  assign rport_io_ins_303 = regOuts_303;
  assign rport_io_ins_304 = regOuts_304;
  assign rport_io_ins_305 = regOuts_305;
  assign rport_io_ins_306 = regOuts_306;
  assign rport_io_ins_307 = regOuts_307;
  assign rport_io_ins_308 = regOuts_308;
  assign rport_io_ins_309 = regOuts_309;
  assign rport_io_ins_310 = regOuts_310;
  assign rport_io_ins_311 = regOuts_311;
  assign rport_io_ins_312 = regOuts_312;
  assign rport_io_ins_313 = regOuts_313;
  assign rport_io_ins_314 = regOuts_314;
  assign rport_io_ins_315 = regOuts_315;
  assign rport_io_ins_316 = regOuts_316;
  assign rport_io_ins_317 = regOuts_317;
  assign rport_io_ins_318 = regOuts_318;
  assign rport_io_ins_319 = regOuts_319;
  assign rport_io_ins_320 = regOuts_320;
  assign rport_io_ins_321 = regOuts_321;
  assign rport_io_ins_322 = regOuts_322;
  assign rport_io_ins_323 = regOuts_323;
  assign rport_io_ins_324 = regOuts_324;
  assign rport_io_ins_325 = regOuts_325;
  assign rport_io_ins_326 = regOuts_326;
  assign rport_io_ins_327 = regOuts_327;
  assign rport_io_ins_328 = regOuts_328;
  assign rport_io_ins_329 = regOuts_329;
  assign rport_io_ins_330 = regOuts_330;
  assign rport_io_ins_331 = regOuts_331;
  assign rport_io_ins_332 = regOuts_332;
  assign rport_io_ins_333 = regOuts_333;
  assign rport_io_ins_334 = regOuts_334;
  assign rport_io_ins_335 = regOuts_335;
  assign rport_io_ins_336 = regOuts_336;
  assign rport_io_ins_337 = regOuts_337;
  assign rport_io_ins_338 = regOuts_338;
  assign rport_io_ins_339 = regOuts_339;
  assign rport_io_ins_340 = regOuts_340;
  assign rport_io_ins_341 = regOuts_341;
  assign rport_io_ins_342 = regOuts_342;
  assign rport_io_ins_343 = regOuts_343;
  assign rport_io_ins_344 = regOuts_344;
  assign rport_io_ins_345 = regOuts_345;
  assign rport_io_ins_346 = regOuts_346;
  assign rport_io_ins_347 = regOuts_347;
  assign rport_io_ins_348 = regOuts_348;
  assign rport_io_ins_349 = regOuts_349;
  assign rport_io_ins_350 = regOuts_350;
  assign rport_io_ins_351 = regOuts_351;
  assign rport_io_ins_352 = regOuts_352;
  assign rport_io_ins_353 = regOuts_353;
  assign rport_io_ins_354 = regOuts_354;
  assign rport_io_ins_355 = regOuts_355;
  assign rport_io_ins_356 = regOuts_356;
  assign rport_io_ins_357 = regOuts_357;
  assign rport_io_ins_358 = regOuts_358;
  assign rport_io_ins_359 = regOuts_359;
  assign rport_io_ins_360 = regOuts_360;
  assign rport_io_ins_361 = regOuts_361;
  assign rport_io_ins_362 = regOuts_362;
  assign rport_io_ins_363 = regOuts_363;
  assign rport_io_ins_364 = regOuts_364;
  assign rport_io_ins_365 = regOuts_365;
  assign rport_io_ins_366 = regOuts_366;
  assign rport_io_ins_367 = regOuts_367;
  assign rport_io_ins_368 = regOuts_368;
  assign rport_io_ins_369 = regOuts_369;
  assign rport_io_ins_370 = regOuts_370;
  assign rport_io_ins_371 = regOuts_371;
  assign rport_io_ins_372 = regOuts_372;
  assign rport_io_ins_373 = regOuts_373;
  assign rport_io_ins_374 = regOuts_374;
  assign rport_io_ins_375 = regOuts_375;
  assign rport_io_ins_376 = regOuts_376;
  assign rport_io_ins_377 = regOuts_377;
  assign rport_io_ins_378 = regOuts_378;
  assign rport_io_ins_379 = regOuts_379;
  assign rport_io_ins_380 = regOuts_380;
  assign rport_io_ins_381 = regOuts_381;
  assign rport_io_ins_382 = regOuts_382;
  assign rport_io_ins_383 = regOuts_383;
  assign rport_io_ins_384 = regOuts_384;
  assign rport_io_ins_385 = regOuts_385;
  assign rport_io_ins_386 = regOuts_386;
  assign rport_io_ins_387 = regOuts_387;
  assign rport_io_ins_388 = regOuts_388;
  assign rport_io_ins_389 = regOuts_389;
  assign rport_io_ins_390 = regOuts_390;
  assign rport_io_ins_391 = regOuts_391;
  assign rport_io_ins_392 = regOuts_392;
  assign rport_io_ins_393 = regOuts_393;
  assign rport_io_ins_394 = regOuts_394;
  assign rport_io_ins_395 = regOuts_395;
  assign rport_io_ins_396 = regOuts_396;
  assign rport_io_ins_397 = regOuts_397;
  assign rport_io_ins_398 = regOuts_398;
  assign rport_io_ins_399 = regOuts_399;
  assign rport_io_ins_400 = regOuts_400;
  assign rport_io_ins_401 = regOuts_401;
  assign rport_io_ins_402 = regOuts_402;
  assign rport_io_ins_403 = regOuts_403;
  assign rport_io_ins_404 = regOuts_404;
  assign rport_io_ins_405 = regOuts_405;
  assign rport_io_ins_406 = regOuts_406;
  assign rport_io_ins_407 = regOuts_407;
  assign rport_io_ins_408 = regOuts_408;
  assign rport_io_ins_409 = regOuts_409;
  assign rport_io_ins_410 = regOuts_410;
  assign rport_io_ins_411 = regOuts_411;
  assign rport_io_ins_412 = regOuts_412;
  assign rport_io_ins_413 = regOuts_413;
  assign rport_io_ins_414 = regOuts_414;
  assign rport_io_ins_415 = regOuts_415;
  assign rport_io_ins_416 = regOuts_416;
  assign rport_io_ins_417 = regOuts_417;
  assign rport_io_ins_418 = regOuts_418;
  assign rport_io_ins_419 = regOuts_419;
  assign rport_io_ins_420 = regOuts_420;
  assign rport_io_ins_421 = regOuts_421;
  assign rport_io_ins_422 = regOuts_422;
  assign rport_io_ins_423 = regOuts_423;
  assign rport_io_ins_424 = regOuts_424;
  assign rport_io_ins_425 = regOuts_425;
  assign rport_io_ins_426 = regOuts_426;
  assign rport_io_ins_427 = regOuts_427;
  assign rport_io_ins_428 = regOuts_428;
  assign rport_io_ins_429 = regOuts_429;
  assign rport_io_ins_430 = regOuts_430;
  assign rport_io_ins_431 = regOuts_431;
  assign rport_io_ins_432 = regOuts_432;
  assign rport_io_ins_433 = regOuts_433;
  assign rport_io_ins_434 = regOuts_434;
  assign rport_io_ins_435 = regOuts_435;
  assign rport_io_ins_436 = regOuts_436;
  assign rport_io_ins_437 = regOuts_437;
  assign rport_io_ins_438 = regOuts_438;
  assign rport_io_ins_439 = regOuts_439;
  assign rport_io_ins_440 = regOuts_440;
  assign rport_io_ins_441 = regOuts_441;
  assign rport_io_ins_442 = regOuts_442;
  assign rport_io_ins_443 = regOuts_443;
  assign rport_io_ins_444 = regOuts_444;
  assign rport_io_ins_445 = regOuts_445;
  assign rport_io_ins_446 = regOuts_446;
  assign rport_io_ins_447 = regOuts_447;
  assign rport_io_ins_448 = regOuts_448;
  assign rport_io_ins_449 = regOuts_449;
  assign rport_io_ins_450 = regOuts_450;
  assign rport_io_ins_451 = regOuts_451;
  assign rport_io_ins_452 = regOuts_452;
  assign rport_io_ins_453 = regOuts_453;
  assign rport_io_ins_454 = regOuts_454;
  assign rport_io_ins_455 = regOuts_455;
  assign rport_io_ins_456 = regOuts_456;
  assign rport_io_ins_457 = regOuts_457;
  assign rport_io_ins_458 = regOuts_458;
  assign rport_io_ins_459 = regOuts_459;
  assign rport_io_ins_460 = regOuts_460;
  assign rport_io_ins_461 = regOuts_461;
  assign rport_io_ins_462 = regOuts_462;
  assign rport_io_ins_463 = regOuts_463;
  assign rport_io_ins_464 = regOuts_464;
  assign rport_io_ins_465 = regOuts_465;
  assign rport_io_ins_466 = regOuts_466;
  assign rport_io_ins_467 = regOuts_467;
  assign rport_io_ins_468 = regOuts_468;
  assign rport_io_ins_469 = regOuts_469;
  assign rport_io_ins_470 = regOuts_470;
  assign rport_io_ins_471 = regOuts_471;
  assign rport_io_ins_472 = regOuts_472;
  assign rport_io_ins_473 = regOuts_473;
  assign rport_io_ins_474 = regOuts_474;
  assign rport_io_ins_475 = regOuts_475;
  assign rport_io_ins_476 = regOuts_476;
  assign rport_io_ins_477 = regOuts_477;
  assign rport_io_ins_478 = regOuts_478;
  assign rport_io_ins_479 = regOuts_479;
  assign rport_io_ins_480 = regOuts_480;
  assign rport_io_ins_481 = regOuts_481;
  assign rport_io_ins_482 = regOuts_482;
  assign rport_io_ins_483 = regOuts_483;
  assign rport_io_ins_484 = regOuts_484;
  assign rport_io_ins_485 = regOuts_485;
  assign rport_io_ins_486 = regOuts_486;
  assign rport_io_ins_487 = regOuts_487;
  assign rport_io_ins_488 = regOuts_488;
  assign rport_io_ins_489 = regOuts_489;
  assign rport_io_ins_490 = regOuts_490;
  assign rport_io_ins_491 = regOuts_491;
  assign rport_io_ins_492 = regOuts_492;
  assign rport_io_ins_493 = regOuts_493;
  assign rport_io_ins_494 = regOuts_494;
  assign rport_io_ins_495 = regOuts_495;
  assign rport_io_ins_496 = regOuts_496;
  assign rport_io_ins_497 = regOuts_497;
  assign rport_io_ins_498 = regOuts_498;
  assign rport_io_ins_499 = regOuts_499;
  assign rport_io_ins_500 = regOuts_500;
  assign rport_io_ins_501 = regOuts_501;
  assign rport_io_ins_502 = regOuts_502;
  assign rport_io_ins_503 = regOuts_503;
  assign rport_io_ins_504 = regOuts_504;
  assign rport_io_sel = io_raddr;
  assign regOuts_0 = regs_0_io_out;
  assign regOuts_1 = regs_1_io_out;
  assign regOuts_2 = regs_2_io_out;
  assign regOuts_3 = regs_3_io_out;
  assign regOuts_4 = regs_4_io_out;
  assign regOuts_5 = regs_5_io_out;
  assign regOuts_6 = regs_6_io_out;
  assign regOuts_7 = regs_7_io_out;
  assign regOuts_8 = regs_8_io_out;
  assign regOuts_9 = regs_9_io_out;
  assign regOuts_10 = regs_10_io_out;
  assign regOuts_11 = regs_11_io_out;
  assign regOuts_12 = regs_12_io_out;
  assign regOuts_13 = regs_13_io_out;
  assign regOuts_14 = regs_14_io_out;
  assign regOuts_15 = regs_15_io_out;
  assign regOuts_16 = regs_16_io_out;
  assign regOuts_17 = regs_17_io_out;
  assign regOuts_18 = regs_18_io_out;
  assign regOuts_19 = regs_19_io_out;
  assign regOuts_20 = regs_20_io_out;
  assign regOuts_21 = regs_21_io_out;
  assign regOuts_22 = regs_22_io_out;
  assign regOuts_23 = regs_23_io_out;
  assign regOuts_24 = regs_24_io_out;
  assign regOuts_25 = regs_25_io_out;
  assign regOuts_26 = regs_26_io_out;
  assign regOuts_27 = regs_27_io_out;
  assign regOuts_28 = regs_28_io_out;
  assign regOuts_29 = regs_29_io_out;
  assign regOuts_30 = regs_30_io_out;
  assign regOuts_31 = regs_31_io_out;
  assign regOuts_32 = regs_32_io_out;
  assign regOuts_33 = regs_33_io_out;
  assign regOuts_34 = regs_34_io_out;
  assign regOuts_35 = regs_35_io_out;
  assign regOuts_36 = regs_36_io_out;
  assign regOuts_37 = regs_37_io_out;
  assign regOuts_38 = regs_38_io_out;
  assign regOuts_39 = regs_39_io_out;
  assign regOuts_40 = regs_40_io_out;
  assign regOuts_41 = regs_41_io_out;
  assign regOuts_42 = regs_42_io_out;
  assign regOuts_43 = regs_43_io_out;
  assign regOuts_44 = regs_44_io_out;
  assign regOuts_45 = regs_45_io_out;
  assign regOuts_46 = regs_46_io_out;
  assign regOuts_47 = regs_47_io_out;
  assign regOuts_48 = regs_48_io_out;
  assign regOuts_49 = regs_49_io_out;
  assign regOuts_50 = regs_50_io_out;
  assign regOuts_51 = regs_51_io_out;
  assign regOuts_52 = regs_52_io_out;
  assign regOuts_53 = regs_53_io_out;
  assign regOuts_54 = regs_54_io_out;
  assign regOuts_55 = regs_55_io_out;
  assign regOuts_56 = regs_56_io_out;
  assign regOuts_57 = regs_57_io_out;
  assign regOuts_58 = regs_58_io_out;
  assign regOuts_59 = regs_59_io_out;
  assign regOuts_60 = regs_60_io_out;
  assign regOuts_61 = regs_61_io_out;
  assign regOuts_62 = regs_62_io_out;
  assign regOuts_63 = regs_63_io_out;
  assign regOuts_64 = regs_64_io_out;
  assign regOuts_65 = regs_65_io_out;
  assign regOuts_66 = regs_66_io_out;
  assign regOuts_67 = regs_67_io_out;
  assign regOuts_68 = regs_68_io_out;
  assign regOuts_69 = regs_69_io_out;
  assign regOuts_70 = regs_70_io_out;
  assign regOuts_71 = regs_71_io_out;
  assign regOuts_72 = regs_72_io_out;
  assign regOuts_73 = regs_73_io_out;
  assign regOuts_74 = regs_74_io_out;
  assign regOuts_75 = regs_75_io_out;
  assign regOuts_76 = regs_76_io_out;
  assign regOuts_77 = regs_77_io_out;
  assign regOuts_78 = regs_78_io_out;
  assign regOuts_79 = regs_79_io_out;
  assign regOuts_80 = regs_80_io_out;
  assign regOuts_81 = regs_81_io_out;
  assign regOuts_82 = regs_82_io_out;
  assign regOuts_83 = regs_83_io_out;
  assign regOuts_84 = regs_84_io_out;
  assign regOuts_85 = regs_85_io_out;
  assign regOuts_86 = regs_86_io_out;
  assign regOuts_87 = regs_87_io_out;
  assign regOuts_88 = regs_88_io_out;
  assign regOuts_89 = regs_89_io_out;
  assign regOuts_90 = regs_90_io_out;
  assign regOuts_91 = regs_91_io_out;
  assign regOuts_92 = regs_92_io_out;
  assign regOuts_93 = regs_93_io_out;
  assign regOuts_94 = regs_94_io_out;
  assign regOuts_95 = regs_95_io_out;
  assign regOuts_96 = regs_96_io_out;
  assign regOuts_97 = regs_97_io_out;
  assign regOuts_98 = regs_98_io_out;
  assign regOuts_99 = regs_99_io_out;
  assign regOuts_100 = regs_100_io_out;
  assign regOuts_101 = regs_101_io_out;
  assign regOuts_102 = regs_102_io_out;
  assign regOuts_103 = regs_103_io_out;
  assign regOuts_104 = regs_104_io_out;
  assign regOuts_105 = regs_105_io_out;
  assign regOuts_106 = regs_106_io_out;
  assign regOuts_107 = regs_107_io_out;
  assign regOuts_108 = regs_108_io_out;
  assign regOuts_109 = regs_109_io_out;
  assign regOuts_110 = regs_110_io_out;
  assign regOuts_111 = regs_111_io_out;
  assign regOuts_112 = regs_112_io_out;
  assign regOuts_113 = regs_113_io_out;
  assign regOuts_114 = regs_114_io_out;
  assign regOuts_115 = regs_115_io_out;
  assign regOuts_116 = regs_116_io_out;
  assign regOuts_117 = regs_117_io_out;
  assign regOuts_118 = regs_118_io_out;
  assign regOuts_119 = regs_119_io_out;
  assign regOuts_120 = regs_120_io_out;
  assign regOuts_121 = regs_121_io_out;
  assign regOuts_122 = regs_122_io_out;
  assign regOuts_123 = regs_123_io_out;
  assign regOuts_124 = regs_124_io_out;
  assign regOuts_125 = regs_125_io_out;
  assign regOuts_126 = regs_126_io_out;
  assign regOuts_127 = regs_127_io_out;
  assign regOuts_128 = regs_128_io_out;
  assign regOuts_129 = regs_129_io_out;
  assign regOuts_130 = regs_130_io_out;
  assign regOuts_131 = regs_131_io_out;
  assign regOuts_132 = regs_132_io_out;
  assign regOuts_133 = regs_133_io_out;
  assign regOuts_134 = regs_134_io_out;
  assign regOuts_135 = regs_135_io_out;
  assign regOuts_136 = regs_136_io_out;
  assign regOuts_137 = regs_137_io_out;
  assign regOuts_138 = regs_138_io_out;
  assign regOuts_139 = regs_139_io_out;
  assign regOuts_140 = regs_140_io_out;
  assign regOuts_141 = regs_141_io_out;
  assign regOuts_142 = regs_142_io_out;
  assign regOuts_143 = regs_143_io_out;
  assign regOuts_144 = regs_144_io_out;
  assign regOuts_145 = regs_145_io_out;
  assign regOuts_146 = regs_146_io_out;
  assign regOuts_147 = regs_147_io_out;
  assign regOuts_148 = regs_148_io_out;
  assign regOuts_149 = regs_149_io_out;
  assign regOuts_150 = regs_150_io_out;
  assign regOuts_151 = regs_151_io_out;
  assign regOuts_152 = regs_152_io_out;
  assign regOuts_153 = regs_153_io_out;
  assign regOuts_154 = regs_154_io_out;
  assign regOuts_155 = regs_155_io_out;
  assign regOuts_156 = regs_156_io_out;
  assign regOuts_157 = regs_157_io_out;
  assign regOuts_158 = regs_158_io_out;
  assign regOuts_159 = regs_159_io_out;
  assign regOuts_160 = regs_160_io_out;
  assign regOuts_161 = regs_161_io_out;
  assign regOuts_162 = regs_162_io_out;
  assign regOuts_163 = regs_163_io_out;
  assign regOuts_164 = regs_164_io_out;
  assign regOuts_165 = regs_165_io_out;
  assign regOuts_166 = regs_166_io_out;
  assign regOuts_167 = regs_167_io_out;
  assign regOuts_168 = regs_168_io_out;
  assign regOuts_169 = regs_169_io_out;
  assign regOuts_170 = regs_170_io_out;
  assign regOuts_171 = regs_171_io_out;
  assign regOuts_172 = regs_172_io_out;
  assign regOuts_173 = regs_173_io_out;
  assign regOuts_174 = regs_174_io_out;
  assign regOuts_175 = regs_175_io_out;
  assign regOuts_176 = regs_176_io_out;
  assign regOuts_177 = regs_177_io_out;
  assign regOuts_178 = regs_178_io_out;
  assign regOuts_179 = regs_179_io_out;
  assign regOuts_180 = regs_180_io_out;
  assign regOuts_181 = regs_181_io_out;
  assign regOuts_182 = regs_182_io_out;
  assign regOuts_183 = regs_183_io_out;
  assign regOuts_184 = regs_184_io_out;
  assign regOuts_185 = regs_185_io_out;
  assign regOuts_186 = regs_186_io_out;
  assign regOuts_187 = regs_187_io_out;
  assign regOuts_188 = regs_188_io_out;
  assign regOuts_189 = regs_189_io_out;
  assign regOuts_190 = regs_190_io_out;
  assign regOuts_191 = regs_191_io_out;
  assign regOuts_192 = regs_192_io_out;
  assign regOuts_193 = regs_193_io_out;
  assign regOuts_194 = regs_194_io_out;
  assign regOuts_195 = regs_195_io_out;
  assign regOuts_196 = regs_196_io_out;
  assign regOuts_197 = regs_197_io_out;
  assign regOuts_198 = regs_198_io_out;
  assign regOuts_199 = regs_199_io_out;
  assign regOuts_200 = regs_200_io_out;
  assign regOuts_201 = regs_201_io_out;
  assign regOuts_202 = regs_202_io_out;
  assign regOuts_203 = regs_203_io_out;
  assign regOuts_204 = regs_204_io_out;
  assign regOuts_205 = regs_205_io_out;
  assign regOuts_206 = regs_206_io_out;
  assign regOuts_207 = regs_207_io_out;
  assign regOuts_208 = regs_208_io_out;
  assign regOuts_209 = regs_209_io_out;
  assign regOuts_210 = regs_210_io_out;
  assign regOuts_211 = regs_211_io_out;
  assign regOuts_212 = regs_212_io_out;
  assign regOuts_213 = regs_213_io_out;
  assign regOuts_214 = regs_214_io_out;
  assign regOuts_215 = regs_215_io_out;
  assign regOuts_216 = regs_216_io_out;
  assign regOuts_217 = regs_217_io_out;
  assign regOuts_218 = regs_218_io_out;
  assign regOuts_219 = regs_219_io_out;
  assign regOuts_220 = regs_220_io_out;
  assign regOuts_221 = regs_221_io_out;
  assign regOuts_222 = regs_222_io_out;
  assign regOuts_223 = regs_223_io_out;
  assign regOuts_224 = regs_224_io_out;
  assign regOuts_225 = regs_225_io_out;
  assign regOuts_226 = regs_226_io_out;
  assign regOuts_227 = regs_227_io_out;
  assign regOuts_228 = regs_228_io_out;
  assign regOuts_229 = regs_229_io_out;
  assign regOuts_230 = regs_230_io_out;
  assign regOuts_231 = regs_231_io_out;
  assign regOuts_232 = regs_232_io_out;
  assign regOuts_233 = regs_233_io_out;
  assign regOuts_234 = regs_234_io_out;
  assign regOuts_235 = regs_235_io_out;
  assign regOuts_236 = regs_236_io_out;
  assign regOuts_237 = regs_237_io_out;
  assign regOuts_238 = regs_238_io_out;
  assign regOuts_239 = regs_239_io_out;
  assign regOuts_240 = regs_240_io_out;
  assign regOuts_241 = regs_241_io_out;
  assign regOuts_242 = regs_242_io_out;
  assign regOuts_243 = regs_243_io_out;
  assign regOuts_244 = regs_244_io_out;
  assign regOuts_245 = regs_245_io_out;
  assign regOuts_246 = regs_246_io_out;
  assign regOuts_247 = regs_247_io_out;
  assign regOuts_248 = regs_248_io_out;
  assign regOuts_249 = regs_249_io_out;
  assign regOuts_250 = regs_250_io_out;
  assign regOuts_251 = regs_251_io_out;
  assign regOuts_252 = regs_252_io_out;
  assign regOuts_253 = regs_253_io_out;
  assign regOuts_254 = regs_254_io_out;
  assign regOuts_255 = regs_255_io_out;
  assign regOuts_256 = regs_256_io_out;
  assign regOuts_257 = regs_257_io_out;
  assign regOuts_258 = regs_258_io_out;
  assign regOuts_259 = regs_259_io_out;
  assign regOuts_260 = regs_260_io_out;
  assign regOuts_261 = regs_261_io_out;
  assign regOuts_262 = regs_262_io_out;
  assign regOuts_263 = regs_263_io_out;
  assign regOuts_264 = regs_264_io_out;
  assign regOuts_265 = regs_265_io_out;
  assign regOuts_266 = regs_266_io_out;
  assign regOuts_267 = regs_267_io_out;
  assign regOuts_268 = regs_268_io_out;
  assign regOuts_269 = regs_269_io_out;
  assign regOuts_270 = regs_270_io_out;
  assign regOuts_271 = regs_271_io_out;
  assign regOuts_272 = regs_272_io_out;
  assign regOuts_273 = regs_273_io_out;
  assign regOuts_274 = regs_274_io_out;
  assign regOuts_275 = regs_275_io_out;
  assign regOuts_276 = regs_276_io_out;
  assign regOuts_277 = regs_277_io_out;
  assign regOuts_278 = regs_278_io_out;
  assign regOuts_279 = regs_279_io_out;
  assign regOuts_280 = regs_280_io_out;
  assign regOuts_281 = regs_281_io_out;
  assign regOuts_282 = regs_282_io_out;
  assign regOuts_283 = regs_283_io_out;
  assign regOuts_284 = regs_284_io_out;
  assign regOuts_285 = regs_285_io_out;
  assign regOuts_286 = regs_286_io_out;
  assign regOuts_287 = regs_287_io_out;
  assign regOuts_288 = regs_288_io_out;
  assign regOuts_289 = regs_289_io_out;
  assign regOuts_290 = regs_290_io_out;
  assign regOuts_291 = regs_291_io_out;
  assign regOuts_292 = regs_292_io_out;
  assign regOuts_293 = regs_293_io_out;
  assign regOuts_294 = regs_294_io_out;
  assign regOuts_295 = regs_295_io_out;
  assign regOuts_296 = regs_296_io_out;
  assign regOuts_297 = regs_297_io_out;
  assign regOuts_298 = regs_298_io_out;
  assign regOuts_299 = regs_299_io_out;
  assign regOuts_300 = regs_300_io_out;
  assign regOuts_301 = regs_301_io_out;
  assign regOuts_302 = regs_302_io_out;
  assign regOuts_303 = regs_303_io_out;
  assign regOuts_304 = regs_304_io_out;
  assign regOuts_305 = regs_305_io_out;
  assign regOuts_306 = regs_306_io_out;
  assign regOuts_307 = regs_307_io_out;
  assign regOuts_308 = regs_308_io_out;
  assign regOuts_309 = regs_309_io_out;
  assign regOuts_310 = regs_310_io_out;
  assign regOuts_311 = regs_311_io_out;
  assign regOuts_312 = regs_312_io_out;
  assign regOuts_313 = regs_313_io_out;
  assign regOuts_314 = regs_314_io_out;
  assign regOuts_315 = regs_315_io_out;
  assign regOuts_316 = regs_316_io_out;
  assign regOuts_317 = regs_317_io_out;
  assign regOuts_318 = regs_318_io_out;
  assign regOuts_319 = regs_319_io_out;
  assign regOuts_320 = regs_320_io_out;
  assign regOuts_321 = regs_321_io_out;
  assign regOuts_322 = regs_322_io_out;
  assign regOuts_323 = regs_323_io_out;
  assign regOuts_324 = regs_324_io_out;
  assign regOuts_325 = regs_325_io_out;
  assign regOuts_326 = regs_326_io_out;
  assign regOuts_327 = regs_327_io_out;
  assign regOuts_328 = regs_328_io_out;
  assign regOuts_329 = regs_329_io_out;
  assign regOuts_330 = regs_330_io_out;
  assign regOuts_331 = regs_331_io_out;
  assign regOuts_332 = regs_332_io_out;
  assign regOuts_333 = regs_333_io_out;
  assign regOuts_334 = regs_334_io_out;
  assign regOuts_335 = regs_335_io_out;
  assign regOuts_336 = regs_336_io_out;
  assign regOuts_337 = regs_337_io_out;
  assign regOuts_338 = regs_338_io_out;
  assign regOuts_339 = regs_339_io_out;
  assign regOuts_340 = regs_340_io_out;
  assign regOuts_341 = regs_341_io_out;
  assign regOuts_342 = regs_342_io_out;
  assign regOuts_343 = regs_343_io_out;
  assign regOuts_344 = regs_344_io_out;
  assign regOuts_345 = regs_345_io_out;
  assign regOuts_346 = regs_346_io_out;
  assign regOuts_347 = regs_347_io_out;
  assign regOuts_348 = regs_348_io_out;
  assign regOuts_349 = regs_349_io_out;
  assign regOuts_350 = regs_350_io_out;
  assign regOuts_351 = regs_351_io_out;
  assign regOuts_352 = regs_352_io_out;
  assign regOuts_353 = regs_353_io_out;
  assign regOuts_354 = regs_354_io_out;
  assign regOuts_355 = regs_355_io_out;
  assign regOuts_356 = regs_356_io_out;
  assign regOuts_357 = regs_357_io_out;
  assign regOuts_358 = regs_358_io_out;
  assign regOuts_359 = regs_359_io_out;
  assign regOuts_360 = regs_360_io_out;
  assign regOuts_361 = regs_361_io_out;
  assign regOuts_362 = regs_362_io_out;
  assign regOuts_363 = regs_363_io_out;
  assign regOuts_364 = regs_364_io_out;
  assign regOuts_365 = regs_365_io_out;
  assign regOuts_366 = regs_366_io_out;
  assign regOuts_367 = regs_367_io_out;
  assign regOuts_368 = regs_368_io_out;
  assign regOuts_369 = regs_369_io_out;
  assign regOuts_370 = regs_370_io_out;
  assign regOuts_371 = regs_371_io_out;
  assign regOuts_372 = regs_372_io_out;
  assign regOuts_373 = regs_373_io_out;
  assign regOuts_374 = regs_374_io_out;
  assign regOuts_375 = regs_375_io_out;
  assign regOuts_376 = regs_376_io_out;
  assign regOuts_377 = regs_377_io_out;
  assign regOuts_378 = regs_378_io_out;
  assign regOuts_379 = regs_379_io_out;
  assign regOuts_380 = regs_380_io_out;
  assign regOuts_381 = regs_381_io_out;
  assign regOuts_382 = regs_382_io_out;
  assign regOuts_383 = regs_383_io_out;
  assign regOuts_384 = regs_384_io_out;
  assign regOuts_385 = regs_385_io_out;
  assign regOuts_386 = regs_386_io_out;
  assign regOuts_387 = regs_387_io_out;
  assign regOuts_388 = regs_388_io_out;
  assign regOuts_389 = regs_389_io_out;
  assign regOuts_390 = regs_390_io_out;
  assign regOuts_391 = regs_391_io_out;
  assign regOuts_392 = regs_392_io_out;
  assign regOuts_393 = regs_393_io_out;
  assign regOuts_394 = regs_394_io_out;
  assign regOuts_395 = regs_395_io_out;
  assign regOuts_396 = regs_396_io_out;
  assign regOuts_397 = regs_397_io_out;
  assign regOuts_398 = regs_398_io_out;
  assign regOuts_399 = regs_399_io_out;
  assign regOuts_400 = regs_400_io_out;
  assign regOuts_401 = regs_401_io_out;
  assign regOuts_402 = regs_402_io_out;
  assign regOuts_403 = regs_403_io_out;
  assign regOuts_404 = regs_404_io_out;
  assign regOuts_405 = regs_405_io_out;
  assign regOuts_406 = regs_406_io_out;
  assign regOuts_407 = regs_407_io_out;
  assign regOuts_408 = regs_408_io_out;
  assign regOuts_409 = regs_409_io_out;
  assign regOuts_410 = regs_410_io_out;
  assign regOuts_411 = regs_411_io_out;
  assign regOuts_412 = regs_412_io_out;
  assign regOuts_413 = regs_413_io_out;
  assign regOuts_414 = regs_414_io_out;
  assign regOuts_415 = regs_415_io_out;
  assign regOuts_416 = regs_416_io_out;
  assign regOuts_417 = regs_417_io_out;
  assign regOuts_418 = regs_418_io_out;
  assign regOuts_419 = regs_419_io_out;
  assign regOuts_420 = regs_420_io_out;
  assign regOuts_421 = regs_421_io_out;
  assign regOuts_422 = regs_422_io_out;
  assign regOuts_423 = regs_423_io_out;
  assign regOuts_424 = regs_424_io_out;
  assign regOuts_425 = regs_425_io_out;
  assign regOuts_426 = regs_426_io_out;
  assign regOuts_427 = regs_427_io_out;
  assign regOuts_428 = regs_428_io_out;
  assign regOuts_429 = regs_429_io_out;
  assign regOuts_430 = regs_430_io_out;
  assign regOuts_431 = regs_431_io_out;
  assign regOuts_432 = regs_432_io_out;
  assign regOuts_433 = regs_433_io_out;
  assign regOuts_434 = regs_434_io_out;
  assign regOuts_435 = regs_435_io_out;
  assign regOuts_436 = regs_436_io_out;
  assign regOuts_437 = regs_437_io_out;
  assign regOuts_438 = regs_438_io_out;
  assign regOuts_439 = regs_439_io_out;
  assign regOuts_440 = regs_440_io_out;
  assign regOuts_441 = regs_441_io_out;
  assign regOuts_442 = regs_442_io_out;
  assign regOuts_443 = regs_443_io_out;
  assign regOuts_444 = regs_444_io_out;
  assign regOuts_445 = regs_445_io_out;
  assign regOuts_446 = regs_446_io_out;
  assign regOuts_447 = regs_447_io_out;
  assign regOuts_448 = regs_448_io_out;
  assign regOuts_449 = regs_449_io_out;
  assign regOuts_450 = regs_450_io_out;
  assign regOuts_451 = regs_451_io_out;
  assign regOuts_452 = regs_452_io_out;
  assign regOuts_453 = regs_453_io_out;
  assign regOuts_454 = regs_454_io_out;
  assign regOuts_455 = regs_455_io_out;
  assign regOuts_456 = regs_456_io_out;
  assign regOuts_457 = regs_457_io_out;
  assign regOuts_458 = regs_458_io_out;
  assign regOuts_459 = regs_459_io_out;
  assign regOuts_460 = regs_460_io_out;
  assign regOuts_461 = regs_461_io_out;
  assign regOuts_462 = regs_462_io_out;
  assign regOuts_463 = regs_463_io_out;
  assign regOuts_464 = regs_464_io_out;
  assign regOuts_465 = regs_465_io_out;
  assign regOuts_466 = regs_466_io_out;
  assign regOuts_467 = regs_467_io_out;
  assign regOuts_468 = regs_468_io_out;
  assign regOuts_469 = regs_469_io_out;
  assign regOuts_470 = regs_470_io_out;
  assign regOuts_471 = regs_471_io_out;
  assign regOuts_472 = regs_472_io_out;
  assign regOuts_473 = regs_473_io_out;
  assign regOuts_474 = regs_474_io_out;
  assign regOuts_475 = regs_475_io_out;
  assign regOuts_476 = regs_476_io_out;
  assign regOuts_477 = regs_477_io_out;
  assign regOuts_478 = regs_478_io_out;
  assign regOuts_479 = regs_479_io_out;
  assign regOuts_480 = regs_480_io_out;
  assign regOuts_481 = regs_481_io_out;
  assign regOuts_482 = regs_482_io_out;
  assign regOuts_483 = regs_483_io_out;
  assign regOuts_484 = regs_484_io_out;
  assign regOuts_485 = regs_485_io_out;
  assign regOuts_486 = regs_486_io_out;
  assign regOuts_487 = regs_487_io_out;
  assign regOuts_488 = regs_488_io_out;
  assign regOuts_489 = regs_489_io_out;
  assign regOuts_490 = regs_490_io_out;
  assign regOuts_491 = regs_491_io_out;
  assign regOuts_492 = regs_492_io_out;
  assign regOuts_493 = regs_493_io_out;
  assign regOuts_494 = regs_494_io_out;
  assign regOuts_495 = regs_495_io_out;
  assign regOuts_496 = regs_496_io_out;
  assign regOuts_497 = regs_497_io_out;
  assign regOuts_498 = regs_498_io_out;
  assign regOuts_499 = regs_499_io_out;
  assign regOuts_500 = regs_500_io_out;
  assign regOuts_501 = regs_501_io_out;
  assign regOuts_502 = regs_502_io_out;
  assign regOuts_503 = regs_503_io_out;
  assign regOuts_504 = regs_504_io_out;
  assign _T_5082_0 = regOuts_0;
  assign _T_5082_1 = regOuts_1;
  assign _T_5082_2 = regOuts_2;
  assign _T_5082_3 = regOuts_3;
endmodule
module RetimeWrapper_675(
  input         clock,
  input         reset,
  input  [39:0] io_in,
  output [39:0] io_out
);
  wire [39:0] sr_out;
  wire [39:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FFType_671(
  input         clock,
  input         reset,
  input  [39:0] io_in,
  output [39:0] io_out,
  input         io_enable
);
  wire [39:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [39:0] RetimeWrapper_io_in;
  wire [39:0] RetimeWrapper_io_out;
  wire [39:0] _T_10;
  wire [39:0] _GEN_0;
  wire [39:0] _GEN_1;
  RetimeWrapper_675 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? 40'h0 : _T_10;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_10;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_10 = RetimeWrapper_io_out;
endmodule
module FF_672(
  input         clock,
  input         reset,
  input  [39:0] io_in,
  output [39:0] io_out,
  input         io_enable
);
  wire  ff_clock;
  wire  ff_reset;
  wire [39:0] ff_io_in;
  wire [39:0] ff_io_out;
  wire  ff_io_enable;
  FFType_671 ff (
    .clock(ff_clock),
    .reset(ff_reset),
    .io_in(ff_io_in),
    .io_out(ff_io_out),
    .io_enable(ff_io_enable)
  );
  assign io_out = ff_io_out;
  assign ff_io_in = io_in;
  assign ff_io_enable = io_enable;
  assign ff_clock = clock;
  assign ff_reset = reset;
endmodule
module Counter_64(
  input   clock,
  input   reset,
  input   io_enable,
  output  io_done
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [39:0] reg$_io_in;
  wire [39:0] reg$_io_out;
  wire  reg$_io_enable;
  wire [40:0] count;
  wire [41:0] _T_12;
  wire [40:0] newval;
  wire  isMax;
  wire [40:0] next;
  wire  _T_14;
  FF_672 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out};
  assign _T_12 = count + 41'h1;
  assign newval = _T_12[40:0];
  assign isMax = newval >= 41'h2cb417800;
  assign next = isMax ? count : newval;
  assign _T_14 = io_enable & isMax;
  assign io_done = _T_14;
  assign reg$_io_in = next[39:0];
  assign reg$_io_enable = io_enable;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module Fringe(
  input         clock,
  input         reset,
  input  [31:0] io_raddr,
  input         io_wen,
  input  [31:0] io_waddr,
  input  [63:0] io_wdata,
  output [63:0] io_rdata,
  output        io_enable,
  input         io_done,
  output [63:0] io_argIns_0,
  output [63:0] io_argIns_1,
  input         io_argOuts_0_valid,
  input  [63:0] io_argOuts_0_bits,
  input         io_dram_0_cmd_ready,
  output        io_dram_0_cmd_valid,
  output [63:0] io_dram_0_cmd_bits_addr,
  output [31:0] io_dram_0_cmd_bits_size,
  output        io_dram_0_cmd_bits_isWr,
  output [25:0] io_dram_0_cmd_bits_tag_uid,
  output [5:0]  io_dram_0_cmd_bits_tag_streamId,
  input         io_dram_0_wdata_ready,
  output        io_dram_0_wdata_valid,
  output [31:0] io_dram_0_wdata_bits_wdata_0,
  output [31:0] io_dram_0_wdata_bits_wdata_1,
  output [31:0] io_dram_0_wdata_bits_wdata_2,
  output [31:0] io_dram_0_wdata_bits_wdata_3,
  output [31:0] io_dram_0_wdata_bits_wdata_4,
  output [31:0] io_dram_0_wdata_bits_wdata_5,
  output [31:0] io_dram_0_wdata_bits_wdata_6,
  output [31:0] io_dram_0_wdata_bits_wdata_7,
  output [31:0] io_dram_0_wdata_bits_wdata_8,
  output [31:0] io_dram_0_wdata_bits_wdata_9,
  output [31:0] io_dram_0_wdata_bits_wdata_10,
  output [31:0] io_dram_0_wdata_bits_wdata_11,
  output [31:0] io_dram_0_wdata_bits_wdata_12,
  output [31:0] io_dram_0_wdata_bits_wdata_13,
  output [31:0] io_dram_0_wdata_bits_wdata_14,
  output [31:0] io_dram_0_wdata_bits_wdata_15,
  output        io_dram_0_wdata_bits_wlast,
  output        io_dram_0_rresp_ready,
  input         io_dram_0_rresp_valid,
  input  [31:0] io_dram_0_rresp_bits_rdata_0,
  input  [31:0] io_dram_0_rresp_bits_rdata_1,
  input  [31:0] io_dram_0_rresp_bits_rdata_2,
  input  [31:0] io_dram_0_rresp_bits_rdata_3,
  input  [31:0] io_dram_0_rresp_bits_rdata_4,
  input  [31:0] io_dram_0_rresp_bits_rdata_5,
  input  [31:0] io_dram_0_rresp_bits_rdata_6,
  input  [31:0] io_dram_0_rresp_bits_rdata_7,
  input  [31:0] io_dram_0_rresp_bits_rdata_8,
  input  [31:0] io_dram_0_rresp_bits_rdata_9,
  input  [31:0] io_dram_0_rresp_bits_rdata_10,
  input  [31:0] io_dram_0_rresp_bits_rdata_11,
  input  [31:0] io_dram_0_rresp_bits_rdata_12,
  input  [31:0] io_dram_0_rresp_bits_rdata_13,
  input  [31:0] io_dram_0_rresp_bits_rdata_14,
  input  [31:0] io_dram_0_rresp_bits_rdata_15,
  input  [5:0]  io_dram_0_rresp_bits_tag_streamId,
  output        io_dram_0_wresp_ready,
  input         io_dram_0_wresp_valid,
  input  [5:0]  io_dram_0_wresp_bits_tag_streamId
);
  wire  mags_0_clock;
  wire  mags_0_reset;
  wire  mags_0_io_enable;
  wire  mags_0_io_dram_cmd_ready;
  wire  mags_0_io_dram_cmd_valid;
  wire [63:0] mags_0_io_dram_cmd_bits_addr;
  wire [31:0] mags_0_io_dram_cmd_bits_size;
  wire  mags_0_io_dram_cmd_bits_isWr;
  wire [25:0] mags_0_io_dram_cmd_bits_tag_uid;
  wire [5:0] mags_0_io_dram_cmd_bits_tag_streamId;
  wire  mags_0_io_dram_wdata_ready;
  wire  mags_0_io_dram_wdata_valid;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_0;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_1;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_2;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_3;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_4;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_5;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_6;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_7;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_8;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_9;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_10;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_11;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_12;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_13;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_14;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_15;
  wire  mags_0_io_dram_wdata_bits_wlast;
  wire  mags_0_io_dram_rresp_ready;
  wire  mags_0_io_dram_rresp_valid;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_0;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_1;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_2;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_3;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_4;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_5;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_6;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_7;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_8;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_9;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_10;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_11;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_12;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_13;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_14;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_15;
  wire [5:0] mags_0_io_dram_rresp_bits_tag_streamId;
  wire  mags_0_io_dram_wresp_ready;
  wire  mags_0_io_dram_wresp_valid;
  wire [5:0] mags_0_io_dram_wresp_bits_tag_streamId;
  wire [31:0] mags_0_io_debugSignals_0;
  wire [31:0] mags_0_io_debugSignals_1;
  wire [31:0] mags_0_io_debugSignals_2;
  wire [31:0] mags_0_io_debugSignals_3;
  wire [31:0] mags_0_io_debugSignals_4;
  wire [31:0] mags_0_io_debugSignals_5;
  wire [31:0] mags_0_io_debugSignals_6;
  wire [31:0] mags_0_io_debugSignals_7;
  wire [31:0] mags_0_io_debugSignals_8;
  wire [31:0] mags_0_io_debugSignals_9;
  wire [31:0] mags_0_io_debugSignals_10;
  wire [31:0] mags_0_io_debugSignals_11;
  wire [31:0] mags_0_io_debugSignals_12;
  wire [31:0] mags_0_io_debugSignals_13;
  wire [31:0] mags_0_io_debugSignals_14;
  wire [31:0] mags_0_io_debugSignals_15;
  wire [31:0] mags_0_io_debugSignals_16;
  wire [31:0] mags_0_io_debugSignals_17;
  wire [31:0] mags_0_io_debugSignals_18;
  wire [31:0] mags_0_io_debugSignals_19;
  wire [31:0] mags_0_io_debugSignals_20;
  wire [31:0] mags_0_io_debugSignals_21;
  wire [31:0] mags_0_io_debugSignals_22;
  wire [31:0] mags_0_io_debugSignals_23;
  wire [31:0] mags_0_io_debugSignals_24;
  wire [31:0] mags_0_io_debugSignals_25;
  wire [31:0] mags_0_io_debugSignals_26;
  wire [31:0] mags_0_io_debugSignals_27;
  wire [31:0] mags_0_io_debugSignals_28;
  wire [31:0] mags_0_io_debugSignals_29;
  wire [31:0] mags_0_io_debugSignals_30;
  wire [31:0] mags_0_io_debugSignals_31;
  wire [31:0] mags_0_io_debugSignals_32;
  wire [31:0] mags_0_io_debugSignals_33;
  wire [31:0] mags_0_io_debugSignals_34;
  wire [31:0] mags_0_io_debugSignals_35;
  wire [31:0] mags_0_io_debugSignals_36;
  wire [31:0] mags_0_io_debugSignals_37;
  wire [31:0] mags_0_io_debugSignals_38;
  wire [31:0] mags_0_io_debugSignals_39;
  wire [31:0] mags_0_io_debugSignals_40;
  wire [31:0] mags_0_io_debugSignals_41;
  wire [31:0] mags_0_io_debugSignals_42;
  wire [31:0] mags_0_io_debugSignals_43;
  wire [31:0] mags_0_io_debugSignals_44;
  wire [31:0] mags_0_io_debugSignals_45;
  wire [31:0] mags_0_io_debugSignals_46;
  wire [31:0] mags_0_io_debugSignals_47;
  wire [31:0] mags_0_io_debugSignals_48;
  wire [31:0] mags_0_io_debugSignals_49;
  wire [31:0] mags_0_io_debugSignals_50;
  wire [31:0] mags_0_io_debugSignals_51;
  wire [31:0] mags_0_io_debugSignals_52;
  wire [31:0] mags_0_io_debugSignals_53;
  wire [31:0] mags_0_io_debugSignals_54;
  wire [31:0] mags_0_io_debugSignals_55;
  wire [31:0] mags_0_io_debugSignals_56;
  wire [31:0] mags_0_io_debugSignals_57;
  wire [31:0] mags_0_io_debugSignals_58;
  wire [31:0] mags_0_io_debugSignals_59;
  wire [31:0] mags_0_io_debugSignals_60;
  wire [31:0] mags_0_io_debugSignals_61;
  wire [31:0] mags_0_io_debugSignals_62;
  wire [31:0] mags_0_io_debugSignals_63;
  wire [31:0] mags_0_io_debugSignals_64;
  wire [31:0] mags_0_io_debugSignals_65;
  wire [31:0] mags_0_io_debugSignals_66;
  wire [31:0] mags_0_io_debugSignals_67;
  wire [31:0] mags_0_io_debugSignals_68;
  wire [31:0] mags_0_io_debugSignals_69;
  wire [31:0] mags_0_io_debugSignals_70;
  wire [31:0] mags_0_io_debugSignals_71;
  wire [31:0] mags_0_io_debugSignals_72;
  wire [31:0] mags_0_io_debugSignals_73;
  wire [31:0] mags_0_io_debugSignals_74;
  wire [31:0] mags_0_io_debugSignals_75;
  wire [31:0] mags_0_io_debugSignals_76;
  wire [31:0] mags_0_io_debugSignals_77;
  wire [31:0] mags_0_io_debugSignals_78;
  wire [31:0] mags_0_io_debugSignals_79;
  wire [31:0] mags_0_io_debugSignals_80;
  wire [31:0] mags_0_io_debugSignals_81;
  wire [31:0] mags_0_io_debugSignals_82;
  wire [31:0] mags_0_io_debugSignals_83;
  wire [31:0] mags_0_io_debugSignals_84;
  wire [31:0] mags_0_io_debugSignals_85;
  wire [31:0] mags_0_io_debugSignals_86;
  wire [31:0] mags_0_io_debugSignals_87;
  wire [31:0] mags_0_io_debugSignals_88;
  wire [31:0] mags_0_io_debugSignals_89;
  wire [31:0] mags_0_io_debugSignals_90;
  wire [31:0] mags_0_io_debugSignals_91;
  wire [31:0] mags_0_io_debugSignals_92;
  wire [31:0] mags_0_io_debugSignals_93;
  wire [31:0] mags_0_io_debugSignals_94;
  wire [31:0] mags_0_io_debugSignals_95;
  wire [31:0] mags_0_io_debugSignals_96;
  wire [31:0] mags_0_io_debugSignals_97;
  wire [31:0] mags_0_io_debugSignals_98;
  wire [31:0] mags_0_io_debugSignals_99;
  wire [31:0] mags_0_io_debugSignals_100;
  wire [31:0] mags_0_io_debugSignals_101;
  wire [31:0] mags_0_io_debugSignals_102;
  wire [31:0] mags_0_io_debugSignals_103;
  wire [31:0] mags_0_io_debugSignals_104;
  wire [31:0] mags_0_io_debugSignals_105;
  wire [31:0] mags_0_io_debugSignals_106;
  wire [31:0] mags_0_io_debugSignals_107;
  wire [31:0] mags_0_io_debugSignals_108;
  wire [31:0] mags_0_io_debugSignals_109;
  wire [31:0] mags_0_io_debugSignals_110;
  wire [31:0] mags_0_io_debugSignals_111;
  wire [31:0] mags_0_io_debugSignals_112;
  wire [31:0] mags_0_io_debugSignals_113;
  wire  regs_clock;
  wire  regs_reset;
  wire [8:0] regs_io_raddr;
  wire  regs_io_wen;
  wire [8:0] regs_io_waddr;
  wire [63:0] regs_io_wdata;
  wire [63:0] regs_io_rdata;
  wire [63:0] regs_io_argIns_0;
  wire [63:0] regs_io_argIns_1;
  wire [63:0] regs_io_argIns_2;
  wire [63:0] regs_io_argIns_3;
  wire  regs_io_argOuts_0_valid;
  wire [63:0] regs_io_argOuts_0_bits;
  wire  regs_io_argOuts_1_valid;
  wire [63:0] regs_io_argOuts_1_bits;
  wire [63:0] regs_io_argOuts_2_bits;
  wire [63:0] regs_io_argOuts_3_bits;
  wire [63:0] regs_io_argOuts_4_bits;
  wire [63:0] regs_io_argOuts_5_bits;
  wire [63:0] regs_io_argOuts_6_bits;
  wire [63:0] regs_io_argOuts_7_bits;
  wire [63:0] regs_io_argOuts_8_bits;
  wire [63:0] regs_io_argOuts_9_bits;
  wire [63:0] regs_io_argOuts_10_bits;
  wire [63:0] regs_io_argOuts_11_bits;
  wire [63:0] regs_io_argOuts_12_bits;
  wire [63:0] regs_io_argOuts_13_bits;
  wire [63:0] regs_io_argOuts_14_bits;
  wire [63:0] regs_io_argOuts_15_bits;
  wire [63:0] regs_io_argOuts_16_bits;
  wire [63:0] regs_io_argOuts_17_bits;
  wire [63:0] regs_io_argOuts_18_bits;
  wire [63:0] regs_io_argOuts_19_bits;
  wire [63:0] regs_io_argOuts_20_bits;
  wire [63:0] regs_io_argOuts_21_bits;
  wire [63:0] regs_io_argOuts_22_bits;
  wire [63:0] regs_io_argOuts_23_bits;
  wire [63:0] regs_io_argOuts_24_bits;
  wire [63:0] regs_io_argOuts_25_bits;
  wire [63:0] regs_io_argOuts_26_bits;
  wire [63:0] regs_io_argOuts_27_bits;
  wire [63:0] regs_io_argOuts_28_bits;
  wire [63:0] regs_io_argOuts_29_bits;
  wire [63:0] regs_io_argOuts_30_bits;
  wire [63:0] regs_io_argOuts_31_bits;
  wire [63:0] regs_io_argOuts_32_bits;
  wire [63:0] regs_io_argOuts_33_bits;
  wire [63:0] regs_io_argOuts_34_bits;
  wire [63:0] regs_io_argOuts_35_bits;
  wire [63:0] regs_io_argOuts_36_bits;
  wire [63:0] regs_io_argOuts_37_bits;
  wire [63:0] regs_io_argOuts_38_bits;
  wire [63:0] regs_io_argOuts_39_bits;
  wire [63:0] regs_io_argOuts_40_bits;
  wire [63:0] regs_io_argOuts_41_bits;
  wire [63:0] regs_io_argOuts_42_bits;
  wire [63:0] regs_io_argOuts_43_bits;
  wire [63:0] regs_io_argOuts_44_bits;
  wire [63:0] regs_io_argOuts_45_bits;
  wire [63:0] regs_io_argOuts_46_bits;
  wire [63:0] regs_io_argOuts_47_bits;
  wire [63:0] regs_io_argOuts_48_bits;
  wire [63:0] regs_io_argOuts_49_bits;
  wire [63:0] regs_io_argOuts_50_bits;
  wire [63:0] regs_io_argOuts_51_bits;
  wire [63:0] regs_io_argOuts_52_bits;
  wire [63:0] regs_io_argOuts_53_bits;
  wire [63:0] regs_io_argOuts_54_bits;
  wire [63:0] regs_io_argOuts_55_bits;
  wire [63:0] regs_io_argOuts_56_bits;
  wire [63:0] regs_io_argOuts_57_bits;
  wire [63:0] regs_io_argOuts_58_bits;
  wire [63:0] regs_io_argOuts_59_bits;
  wire [63:0] regs_io_argOuts_60_bits;
  wire [63:0] regs_io_argOuts_61_bits;
  wire [63:0] regs_io_argOuts_62_bits;
  wire [63:0] regs_io_argOuts_63_bits;
  wire [63:0] regs_io_argOuts_64_bits;
  wire [63:0] regs_io_argOuts_65_bits;
  wire [63:0] regs_io_argOuts_66_bits;
  wire [63:0] regs_io_argOuts_67_bits;
  wire [63:0] regs_io_argOuts_68_bits;
  wire [63:0] regs_io_argOuts_69_bits;
  wire [63:0] regs_io_argOuts_70_bits;
  wire [63:0] regs_io_argOuts_71_bits;
  wire [63:0] regs_io_argOuts_72_bits;
  wire [63:0] regs_io_argOuts_73_bits;
  wire [63:0] regs_io_argOuts_74_bits;
  wire [63:0] regs_io_argOuts_75_bits;
  wire [63:0] regs_io_argOuts_76_bits;
  wire [63:0] regs_io_argOuts_77_bits;
  wire [63:0] regs_io_argOuts_78_bits;
  wire [63:0] regs_io_argOuts_79_bits;
  wire [63:0] regs_io_argOuts_80_bits;
  wire [63:0] regs_io_argOuts_81_bits;
  wire [63:0] regs_io_argOuts_82_bits;
  wire [63:0] regs_io_argOuts_83_bits;
  wire [63:0] regs_io_argOuts_84_bits;
  wire [63:0] regs_io_argOuts_85_bits;
  wire [63:0] regs_io_argOuts_86_bits;
  wire [63:0] regs_io_argOuts_87_bits;
  wire [63:0] regs_io_argOuts_88_bits;
  wire [63:0] regs_io_argOuts_89_bits;
  wire [63:0] regs_io_argOuts_90_bits;
  wire [63:0] regs_io_argOuts_91_bits;
  wire [63:0] regs_io_argOuts_92_bits;
  wire [63:0] regs_io_argOuts_93_bits;
  wire [63:0] regs_io_argOuts_94_bits;
  wire [63:0] regs_io_argOuts_95_bits;
  wire [63:0] regs_io_argOuts_96_bits;
  wire [63:0] regs_io_argOuts_97_bits;
  wire [63:0] regs_io_argOuts_98_bits;
  wire [63:0] regs_io_argOuts_99_bits;
  wire [63:0] regs_io_argOuts_100_bits;
  wire [63:0] regs_io_argOuts_101_bits;
  wire [63:0] regs_io_argOuts_102_bits;
  wire [63:0] regs_io_argOuts_103_bits;
  wire [63:0] regs_io_argOuts_104_bits;
  wire [63:0] regs_io_argOuts_105_bits;
  wire [63:0] regs_io_argOuts_106_bits;
  wire [63:0] regs_io_argOuts_107_bits;
  wire [63:0] regs_io_argOuts_108_bits;
  wire [63:0] regs_io_argOuts_109_bits;
  wire [63:0] regs_io_argOuts_110_bits;
  wire [63:0] regs_io_argOuts_111_bits;
  wire [63:0] regs_io_argOuts_112_bits;
  wire [63:0] regs_io_argOuts_113_bits;
  wire [63:0] regs_io_argOuts_114_bits;
  wire [63:0] regs_io_argOuts_115_bits;
  reg [63:0] _T_524;
  reg [63:0] _RAND_0;
  wire [63:0] _GEN_0;
  wire  _T_525;
  wire  _T_526;
  wire  _T_527;
  wire  localEnable;
  wire  timeoutCtr_clock;
  wire  timeoutCtr_reset;
  wire  timeoutCtr_io_enable;
  wire  timeoutCtr_io_done;
  wire  depulser_clock;
  wire  depulser_reset;
  wire  depulser_io_in;
  wire  depulser_io_rst;
  wire  depulser_io_out;
  wire  _T_532;
  wire [63:0] _T_533;
  wire  status_valid;
  wire [63:0] status_bits;
  wire  _T_543;
  wire  _T_545;
  wire [1:0] _T_546;
  MAGCore mags_0 (
    .clock(mags_0_clock),
    .reset(mags_0_reset),
    .io_enable(mags_0_io_enable),
    .io_dram_cmd_ready(mags_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(mags_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(mags_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(mags_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(mags_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag_uid(mags_0_io_dram_cmd_bits_tag_uid),
    .io_dram_cmd_bits_tag_streamId(mags_0_io_dram_cmd_bits_tag_streamId),
    .io_dram_wdata_ready(mags_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(mags_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(mags_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(mags_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(mags_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(mags_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(mags_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(mags_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(mags_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(mags_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(mags_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(mags_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(mags_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(mags_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(mags_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(mags_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(mags_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(mags_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wlast(mags_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(mags_0_io_dram_rresp_ready),
    .io_dram_rresp_valid(mags_0_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(mags_0_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(mags_0_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(mags_0_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(mags_0_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(mags_0_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(mags_0_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(mags_0_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(mags_0_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_rdata_8(mags_0_io_dram_rresp_bits_rdata_8),
    .io_dram_rresp_bits_rdata_9(mags_0_io_dram_rresp_bits_rdata_9),
    .io_dram_rresp_bits_rdata_10(mags_0_io_dram_rresp_bits_rdata_10),
    .io_dram_rresp_bits_rdata_11(mags_0_io_dram_rresp_bits_rdata_11),
    .io_dram_rresp_bits_rdata_12(mags_0_io_dram_rresp_bits_rdata_12),
    .io_dram_rresp_bits_rdata_13(mags_0_io_dram_rresp_bits_rdata_13),
    .io_dram_rresp_bits_rdata_14(mags_0_io_dram_rresp_bits_rdata_14),
    .io_dram_rresp_bits_rdata_15(mags_0_io_dram_rresp_bits_rdata_15),
    .io_dram_rresp_bits_tag_streamId(mags_0_io_dram_rresp_bits_tag_streamId),
    .io_dram_wresp_ready(mags_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(mags_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag_streamId(mags_0_io_dram_wresp_bits_tag_streamId),
    .io_debugSignals_0(mags_0_io_debugSignals_0),
    .io_debugSignals_1(mags_0_io_debugSignals_1),
    .io_debugSignals_2(mags_0_io_debugSignals_2),
    .io_debugSignals_3(mags_0_io_debugSignals_3),
    .io_debugSignals_4(mags_0_io_debugSignals_4),
    .io_debugSignals_5(mags_0_io_debugSignals_5),
    .io_debugSignals_6(mags_0_io_debugSignals_6),
    .io_debugSignals_7(mags_0_io_debugSignals_7),
    .io_debugSignals_8(mags_0_io_debugSignals_8),
    .io_debugSignals_9(mags_0_io_debugSignals_9),
    .io_debugSignals_10(mags_0_io_debugSignals_10),
    .io_debugSignals_11(mags_0_io_debugSignals_11),
    .io_debugSignals_12(mags_0_io_debugSignals_12),
    .io_debugSignals_13(mags_0_io_debugSignals_13),
    .io_debugSignals_14(mags_0_io_debugSignals_14),
    .io_debugSignals_15(mags_0_io_debugSignals_15),
    .io_debugSignals_16(mags_0_io_debugSignals_16),
    .io_debugSignals_17(mags_0_io_debugSignals_17),
    .io_debugSignals_18(mags_0_io_debugSignals_18),
    .io_debugSignals_19(mags_0_io_debugSignals_19),
    .io_debugSignals_20(mags_0_io_debugSignals_20),
    .io_debugSignals_21(mags_0_io_debugSignals_21),
    .io_debugSignals_22(mags_0_io_debugSignals_22),
    .io_debugSignals_23(mags_0_io_debugSignals_23),
    .io_debugSignals_24(mags_0_io_debugSignals_24),
    .io_debugSignals_25(mags_0_io_debugSignals_25),
    .io_debugSignals_26(mags_0_io_debugSignals_26),
    .io_debugSignals_27(mags_0_io_debugSignals_27),
    .io_debugSignals_28(mags_0_io_debugSignals_28),
    .io_debugSignals_29(mags_0_io_debugSignals_29),
    .io_debugSignals_30(mags_0_io_debugSignals_30),
    .io_debugSignals_31(mags_0_io_debugSignals_31),
    .io_debugSignals_32(mags_0_io_debugSignals_32),
    .io_debugSignals_33(mags_0_io_debugSignals_33),
    .io_debugSignals_34(mags_0_io_debugSignals_34),
    .io_debugSignals_35(mags_0_io_debugSignals_35),
    .io_debugSignals_36(mags_0_io_debugSignals_36),
    .io_debugSignals_37(mags_0_io_debugSignals_37),
    .io_debugSignals_38(mags_0_io_debugSignals_38),
    .io_debugSignals_39(mags_0_io_debugSignals_39),
    .io_debugSignals_40(mags_0_io_debugSignals_40),
    .io_debugSignals_41(mags_0_io_debugSignals_41),
    .io_debugSignals_42(mags_0_io_debugSignals_42),
    .io_debugSignals_43(mags_0_io_debugSignals_43),
    .io_debugSignals_44(mags_0_io_debugSignals_44),
    .io_debugSignals_45(mags_0_io_debugSignals_45),
    .io_debugSignals_46(mags_0_io_debugSignals_46),
    .io_debugSignals_47(mags_0_io_debugSignals_47),
    .io_debugSignals_48(mags_0_io_debugSignals_48),
    .io_debugSignals_49(mags_0_io_debugSignals_49),
    .io_debugSignals_50(mags_0_io_debugSignals_50),
    .io_debugSignals_51(mags_0_io_debugSignals_51),
    .io_debugSignals_52(mags_0_io_debugSignals_52),
    .io_debugSignals_53(mags_0_io_debugSignals_53),
    .io_debugSignals_54(mags_0_io_debugSignals_54),
    .io_debugSignals_55(mags_0_io_debugSignals_55),
    .io_debugSignals_56(mags_0_io_debugSignals_56),
    .io_debugSignals_57(mags_0_io_debugSignals_57),
    .io_debugSignals_58(mags_0_io_debugSignals_58),
    .io_debugSignals_59(mags_0_io_debugSignals_59),
    .io_debugSignals_60(mags_0_io_debugSignals_60),
    .io_debugSignals_61(mags_0_io_debugSignals_61),
    .io_debugSignals_62(mags_0_io_debugSignals_62),
    .io_debugSignals_63(mags_0_io_debugSignals_63),
    .io_debugSignals_64(mags_0_io_debugSignals_64),
    .io_debugSignals_65(mags_0_io_debugSignals_65),
    .io_debugSignals_66(mags_0_io_debugSignals_66),
    .io_debugSignals_67(mags_0_io_debugSignals_67),
    .io_debugSignals_68(mags_0_io_debugSignals_68),
    .io_debugSignals_69(mags_0_io_debugSignals_69),
    .io_debugSignals_70(mags_0_io_debugSignals_70),
    .io_debugSignals_71(mags_0_io_debugSignals_71),
    .io_debugSignals_72(mags_0_io_debugSignals_72),
    .io_debugSignals_73(mags_0_io_debugSignals_73),
    .io_debugSignals_74(mags_0_io_debugSignals_74),
    .io_debugSignals_75(mags_0_io_debugSignals_75),
    .io_debugSignals_76(mags_0_io_debugSignals_76),
    .io_debugSignals_77(mags_0_io_debugSignals_77),
    .io_debugSignals_78(mags_0_io_debugSignals_78),
    .io_debugSignals_79(mags_0_io_debugSignals_79),
    .io_debugSignals_80(mags_0_io_debugSignals_80),
    .io_debugSignals_81(mags_0_io_debugSignals_81),
    .io_debugSignals_82(mags_0_io_debugSignals_82),
    .io_debugSignals_83(mags_0_io_debugSignals_83),
    .io_debugSignals_84(mags_0_io_debugSignals_84),
    .io_debugSignals_85(mags_0_io_debugSignals_85),
    .io_debugSignals_86(mags_0_io_debugSignals_86),
    .io_debugSignals_87(mags_0_io_debugSignals_87),
    .io_debugSignals_88(mags_0_io_debugSignals_88),
    .io_debugSignals_89(mags_0_io_debugSignals_89),
    .io_debugSignals_90(mags_0_io_debugSignals_90),
    .io_debugSignals_91(mags_0_io_debugSignals_91),
    .io_debugSignals_92(mags_0_io_debugSignals_92),
    .io_debugSignals_93(mags_0_io_debugSignals_93),
    .io_debugSignals_94(mags_0_io_debugSignals_94),
    .io_debugSignals_95(mags_0_io_debugSignals_95),
    .io_debugSignals_96(mags_0_io_debugSignals_96),
    .io_debugSignals_97(mags_0_io_debugSignals_97),
    .io_debugSignals_98(mags_0_io_debugSignals_98),
    .io_debugSignals_99(mags_0_io_debugSignals_99),
    .io_debugSignals_100(mags_0_io_debugSignals_100),
    .io_debugSignals_101(mags_0_io_debugSignals_101),
    .io_debugSignals_102(mags_0_io_debugSignals_102),
    .io_debugSignals_103(mags_0_io_debugSignals_103),
    .io_debugSignals_104(mags_0_io_debugSignals_104),
    .io_debugSignals_105(mags_0_io_debugSignals_105),
    .io_debugSignals_106(mags_0_io_debugSignals_106),
    .io_debugSignals_107(mags_0_io_debugSignals_107),
    .io_debugSignals_108(mags_0_io_debugSignals_108),
    .io_debugSignals_109(mags_0_io_debugSignals_109),
    .io_debugSignals_110(mags_0_io_debugSignals_110),
    .io_debugSignals_111(mags_0_io_debugSignals_111),
    .io_debugSignals_112(mags_0_io_debugSignals_112),
    .io_debugSignals_113(mags_0_io_debugSignals_113)
  );
  RegFile regs (
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits),
    .io_argOuts_2_bits(regs_io_argOuts_2_bits),
    .io_argOuts_3_bits(regs_io_argOuts_3_bits),
    .io_argOuts_4_bits(regs_io_argOuts_4_bits),
    .io_argOuts_5_bits(regs_io_argOuts_5_bits),
    .io_argOuts_6_bits(regs_io_argOuts_6_bits),
    .io_argOuts_7_bits(regs_io_argOuts_7_bits),
    .io_argOuts_8_bits(regs_io_argOuts_8_bits),
    .io_argOuts_9_bits(regs_io_argOuts_9_bits),
    .io_argOuts_10_bits(regs_io_argOuts_10_bits),
    .io_argOuts_11_bits(regs_io_argOuts_11_bits),
    .io_argOuts_12_bits(regs_io_argOuts_12_bits),
    .io_argOuts_13_bits(regs_io_argOuts_13_bits),
    .io_argOuts_14_bits(regs_io_argOuts_14_bits),
    .io_argOuts_15_bits(regs_io_argOuts_15_bits),
    .io_argOuts_16_bits(regs_io_argOuts_16_bits),
    .io_argOuts_17_bits(regs_io_argOuts_17_bits),
    .io_argOuts_18_bits(regs_io_argOuts_18_bits),
    .io_argOuts_19_bits(regs_io_argOuts_19_bits),
    .io_argOuts_20_bits(regs_io_argOuts_20_bits),
    .io_argOuts_21_bits(regs_io_argOuts_21_bits),
    .io_argOuts_22_bits(regs_io_argOuts_22_bits),
    .io_argOuts_23_bits(regs_io_argOuts_23_bits),
    .io_argOuts_24_bits(regs_io_argOuts_24_bits),
    .io_argOuts_25_bits(regs_io_argOuts_25_bits),
    .io_argOuts_26_bits(regs_io_argOuts_26_bits),
    .io_argOuts_27_bits(regs_io_argOuts_27_bits),
    .io_argOuts_28_bits(regs_io_argOuts_28_bits),
    .io_argOuts_29_bits(regs_io_argOuts_29_bits),
    .io_argOuts_30_bits(regs_io_argOuts_30_bits),
    .io_argOuts_31_bits(regs_io_argOuts_31_bits),
    .io_argOuts_32_bits(regs_io_argOuts_32_bits),
    .io_argOuts_33_bits(regs_io_argOuts_33_bits),
    .io_argOuts_34_bits(regs_io_argOuts_34_bits),
    .io_argOuts_35_bits(regs_io_argOuts_35_bits),
    .io_argOuts_36_bits(regs_io_argOuts_36_bits),
    .io_argOuts_37_bits(regs_io_argOuts_37_bits),
    .io_argOuts_38_bits(regs_io_argOuts_38_bits),
    .io_argOuts_39_bits(regs_io_argOuts_39_bits),
    .io_argOuts_40_bits(regs_io_argOuts_40_bits),
    .io_argOuts_41_bits(regs_io_argOuts_41_bits),
    .io_argOuts_42_bits(regs_io_argOuts_42_bits),
    .io_argOuts_43_bits(regs_io_argOuts_43_bits),
    .io_argOuts_44_bits(regs_io_argOuts_44_bits),
    .io_argOuts_45_bits(regs_io_argOuts_45_bits),
    .io_argOuts_46_bits(regs_io_argOuts_46_bits),
    .io_argOuts_47_bits(regs_io_argOuts_47_bits),
    .io_argOuts_48_bits(regs_io_argOuts_48_bits),
    .io_argOuts_49_bits(regs_io_argOuts_49_bits),
    .io_argOuts_50_bits(regs_io_argOuts_50_bits),
    .io_argOuts_51_bits(regs_io_argOuts_51_bits),
    .io_argOuts_52_bits(regs_io_argOuts_52_bits),
    .io_argOuts_53_bits(regs_io_argOuts_53_bits),
    .io_argOuts_54_bits(regs_io_argOuts_54_bits),
    .io_argOuts_55_bits(regs_io_argOuts_55_bits),
    .io_argOuts_56_bits(regs_io_argOuts_56_bits),
    .io_argOuts_57_bits(regs_io_argOuts_57_bits),
    .io_argOuts_58_bits(regs_io_argOuts_58_bits),
    .io_argOuts_59_bits(regs_io_argOuts_59_bits),
    .io_argOuts_60_bits(regs_io_argOuts_60_bits),
    .io_argOuts_61_bits(regs_io_argOuts_61_bits),
    .io_argOuts_62_bits(regs_io_argOuts_62_bits),
    .io_argOuts_63_bits(regs_io_argOuts_63_bits),
    .io_argOuts_64_bits(regs_io_argOuts_64_bits),
    .io_argOuts_65_bits(regs_io_argOuts_65_bits),
    .io_argOuts_66_bits(regs_io_argOuts_66_bits),
    .io_argOuts_67_bits(regs_io_argOuts_67_bits),
    .io_argOuts_68_bits(regs_io_argOuts_68_bits),
    .io_argOuts_69_bits(regs_io_argOuts_69_bits),
    .io_argOuts_70_bits(regs_io_argOuts_70_bits),
    .io_argOuts_71_bits(regs_io_argOuts_71_bits),
    .io_argOuts_72_bits(regs_io_argOuts_72_bits),
    .io_argOuts_73_bits(regs_io_argOuts_73_bits),
    .io_argOuts_74_bits(regs_io_argOuts_74_bits),
    .io_argOuts_75_bits(regs_io_argOuts_75_bits),
    .io_argOuts_76_bits(regs_io_argOuts_76_bits),
    .io_argOuts_77_bits(regs_io_argOuts_77_bits),
    .io_argOuts_78_bits(regs_io_argOuts_78_bits),
    .io_argOuts_79_bits(regs_io_argOuts_79_bits),
    .io_argOuts_80_bits(regs_io_argOuts_80_bits),
    .io_argOuts_81_bits(regs_io_argOuts_81_bits),
    .io_argOuts_82_bits(regs_io_argOuts_82_bits),
    .io_argOuts_83_bits(regs_io_argOuts_83_bits),
    .io_argOuts_84_bits(regs_io_argOuts_84_bits),
    .io_argOuts_85_bits(regs_io_argOuts_85_bits),
    .io_argOuts_86_bits(regs_io_argOuts_86_bits),
    .io_argOuts_87_bits(regs_io_argOuts_87_bits),
    .io_argOuts_88_bits(regs_io_argOuts_88_bits),
    .io_argOuts_89_bits(regs_io_argOuts_89_bits),
    .io_argOuts_90_bits(regs_io_argOuts_90_bits),
    .io_argOuts_91_bits(regs_io_argOuts_91_bits),
    .io_argOuts_92_bits(regs_io_argOuts_92_bits),
    .io_argOuts_93_bits(regs_io_argOuts_93_bits),
    .io_argOuts_94_bits(regs_io_argOuts_94_bits),
    .io_argOuts_95_bits(regs_io_argOuts_95_bits),
    .io_argOuts_96_bits(regs_io_argOuts_96_bits),
    .io_argOuts_97_bits(regs_io_argOuts_97_bits),
    .io_argOuts_98_bits(regs_io_argOuts_98_bits),
    .io_argOuts_99_bits(regs_io_argOuts_99_bits),
    .io_argOuts_100_bits(regs_io_argOuts_100_bits),
    .io_argOuts_101_bits(regs_io_argOuts_101_bits),
    .io_argOuts_102_bits(regs_io_argOuts_102_bits),
    .io_argOuts_103_bits(regs_io_argOuts_103_bits),
    .io_argOuts_104_bits(regs_io_argOuts_104_bits),
    .io_argOuts_105_bits(regs_io_argOuts_105_bits),
    .io_argOuts_106_bits(regs_io_argOuts_106_bits),
    .io_argOuts_107_bits(regs_io_argOuts_107_bits),
    .io_argOuts_108_bits(regs_io_argOuts_108_bits),
    .io_argOuts_109_bits(regs_io_argOuts_109_bits),
    .io_argOuts_110_bits(regs_io_argOuts_110_bits),
    .io_argOuts_111_bits(regs_io_argOuts_111_bits),
    .io_argOuts_112_bits(regs_io_argOuts_112_bits),
    .io_argOuts_113_bits(regs_io_argOuts_113_bits),
    .io_argOuts_114_bits(regs_io_argOuts_114_bits),
    .io_argOuts_115_bits(regs_io_argOuts_115_bits)
  );
  Counter_64 timeoutCtr (
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser (
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _GEN_0 = regs_io_rdata;
  assign _T_525 = regs_io_argIns_0[0];
  assign _T_526 = regs_io_argIns_1[0];
  assign _T_527 = ~ _T_526;
  assign localEnable = _T_525 & _T_527;
  assign _T_532 = io_done | timeoutCtr_io_done;
  assign _T_533 = ~ regs_io_argIns_0;
  assign _T_543 = _T_525 & timeoutCtr_io_done;
  assign _T_545 = _T_525 & depulser_io_out;
  assign _T_546 = {_T_543,_T_545};
  assign io_rdata = _T_524;
  assign io_enable = localEnable;
  assign io_argIns_0 = regs_io_argIns_2;
  assign io_argIns_1 = regs_io_argIns_3;
  assign io_dram_0_cmd_valid = mags_0_io_dram_cmd_valid;
  assign io_dram_0_cmd_bits_addr = mags_0_io_dram_cmd_bits_addr;
  assign io_dram_0_cmd_bits_size = mags_0_io_dram_cmd_bits_size;
  assign io_dram_0_cmd_bits_isWr = mags_0_io_dram_cmd_bits_isWr;
  assign io_dram_0_cmd_bits_tag_uid = mags_0_io_dram_cmd_bits_tag_uid;
  assign io_dram_0_cmd_bits_tag_streamId = mags_0_io_dram_cmd_bits_tag_streamId;
  assign io_dram_0_wdata_valid = mags_0_io_dram_wdata_valid;
  assign io_dram_0_wdata_bits_wdata_0 = mags_0_io_dram_wdata_bits_wdata_0;
  assign io_dram_0_wdata_bits_wdata_1 = mags_0_io_dram_wdata_bits_wdata_1;
  assign io_dram_0_wdata_bits_wdata_2 = mags_0_io_dram_wdata_bits_wdata_2;
  assign io_dram_0_wdata_bits_wdata_3 = mags_0_io_dram_wdata_bits_wdata_3;
  assign io_dram_0_wdata_bits_wdata_4 = mags_0_io_dram_wdata_bits_wdata_4;
  assign io_dram_0_wdata_bits_wdata_5 = mags_0_io_dram_wdata_bits_wdata_5;
  assign io_dram_0_wdata_bits_wdata_6 = mags_0_io_dram_wdata_bits_wdata_6;
  assign io_dram_0_wdata_bits_wdata_7 = mags_0_io_dram_wdata_bits_wdata_7;
  assign io_dram_0_wdata_bits_wdata_8 = mags_0_io_dram_wdata_bits_wdata_8;
  assign io_dram_0_wdata_bits_wdata_9 = mags_0_io_dram_wdata_bits_wdata_9;
  assign io_dram_0_wdata_bits_wdata_10 = mags_0_io_dram_wdata_bits_wdata_10;
  assign io_dram_0_wdata_bits_wdata_11 = mags_0_io_dram_wdata_bits_wdata_11;
  assign io_dram_0_wdata_bits_wdata_12 = mags_0_io_dram_wdata_bits_wdata_12;
  assign io_dram_0_wdata_bits_wdata_13 = mags_0_io_dram_wdata_bits_wdata_13;
  assign io_dram_0_wdata_bits_wdata_14 = mags_0_io_dram_wdata_bits_wdata_14;
  assign io_dram_0_wdata_bits_wdata_15 = mags_0_io_dram_wdata_bits_wdata_15;
  assign io_dram_0_wdata_bits_wlast = mags_0_io_dram_wdata_bits_wlast;
  assign io_dram_0_rresp_ready = mags_0_io_dram_rresp_ready;
  assign io_dram_0_wresp_ready = mags_0_io_dram_wresp_ready;
  assign mags_0_io_enable = localEnable;
  assign mags_0_io_dram_cmd_ready = io_dram_0_cmd_ready;
  assign mags_0_io_dram_wdata_ready = io_dram_0_wdata_ready;
  assign mags_0_io_dram_rresp_valid = io_dram_0_rresp_valid;
  assign mags_0_io_dram_rresp_bits_rdata_0 = io_dram_0_rresp_bits_rdata_0;
  assign mags_0_io_dram_rresp_bits_rdata_1 = io_dram_0_rresp_bits_rdata_1;
  assign mags_0_io_dram_rresp_bits_rdata_2 = io_dram_0_rresp_bits_rdata_2;
  assign mags_0_io_dram_rresp_bits_rdata_3 = io_dram_0_rresp_bits_rdata_3;
  assign mags_0_io_dram_rresp_bits_rdata_4 = io_dram_0_rresp_bits_rdata_4;
  assign mags_0_io_dram_rresp_bits_rdata_5 = io_dram_0_rresp_bits_rdata_5;
  assign mags_0_io_dram_rresp_bits_rdata_6 = io_dram_0_rresp_bits_rdata_6;
  assign mags_0_io_dram_rresp_bits_rdata_7 = io_dram_0_rresp_bits_rdata_7;
  assign mags_0_io_dram_rresp_bits_rdata_8 = io_dram_0_rresp_bits_rdata_8;
  assign mags_0_io_dram_rresp_bits_rdata_9 = io_dram_0_rresp_bits_rdata_9;
  assign mags_0_io_dram_rresp_bits_rdata_10 = io_dram_0_rresp_bits_rdata_10;
  assign mags_0_io_dram_rresp_bits_rdata_11 = io_dram_0_rresp_bits_rdata_11;
  assign mags_0_io_dram_rresp_bits_rdata_12 = io_dram_0_rresp_bits_rdata_12;
  assign mags_0_io_dram_rresp_bits_rdata_13 = io_dram_0_rresp_bits_rdata_13;
  assign mags_0_io_dram_rresp_bits_rdata_14 = io_dram_0_rresp_bits_rdata_14;
  assign mags_0_io_dram_rresp_bits_rdata_15 = io_dram_0_rresp_bits_rdata_15;
  assign mags_0_io_dram_rresp_bits_tag_streamId = io_dram_0_rresp_bits_tag_streamId;
  assign mags_0_io_dram_wresp_valid = io_dram_0_wresp_valid;
  assign mags_0_io_dram_wresp_bits_tag_streamId = io_dram_0_wresp_bits_tag_streamId;
  assign mags_0_clock = clock;
  assign mags_0_reset = reset;
  assign regs_io_raddr = io_raddr[8:0];
  assign regs_io_wen = io_wen;
  assign regs_io_waddr = io_waddr[8:0];
  assign regs_io_wdata = io_wdata;
  assign regs_io_argOuts_0_valid = status_valid;
  assign regs_io_argOuts_0_bits = status_bits;
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid;
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits;
  assign regs_io_argOuts_2_bits = {{32'd0}, mags_0_io_debugSignals_0};
  assign regs_io_argOuts_3_bits = {{32'd0}, mags_0_io_debugSignals_1};
  assign regs_io_argOuts_4_bits = {{32'd0}, mags_0_io_debugSignals_2};
  assign regs_io_argOuts_5_bits = {{32'd0}, mags_0_io_debugSignals_3};
  assign regs_io_argOuts_6_bits = {{32'd0}, mags_0_io_debugSignals_4};
  assign regs_io_argOuts_7_bits = {{32'd0}, mags_0_io_debugSignals_5};
  assign regs_io_argOuts_8_bits = {{32'd0}, mags_0_io_debugSignals_6};
  assign regs_io_argOuts_9_bits = {{32'd0}, mags_0_io_debugSignals_7};
  assign regs_io_argOuts_10_bits = {{32'd0}, mags_0_io_debugSignals_8};
  assign regs_io_argOuts_11_bits = {{32'd0}, mags_0_io_debugSignals_9};
  assign regs_io_argOuts_12_bits = {{32'd0}, mags_0_io_debugSignals_10};
  assign regs_io_argOuts_13_bits = {{32'd0}, mags_0_io_debugSignals_11};
  assign regs_io_argOuts_14_bits = {{32'd0}, mags_0_io_debugSignals_12};
  assign regs_io_argOuts_15_bits = {{32'd0}, mags_0_io_debugSignals_13};
  assign regs_io_argOuts_16_bits = {{32'd0}, mags_0_io_debugSignals_14};
  assign regs_io_argOuts_17_bits = {{32'd0}, mags_0_io_debugSignals_15};
  assign regs_io_argOuts_18_bits = {{32'd0}, mags_0_io_debugSignals_16};
  assign regs_io_argOuts_19_bits = {{32'd0}, mags_0_io_debugSignals_17};
  assign regs_io_argOuts_20_bits = {{32'd0}, mags_0_io_debugSignals_18};
  assign regs_io_argOuts_21_bits = {{32'd0}, mags_0_io_debugSignals_19};
  assign regs_io_argOuts_22_bits = {{32'd0}, mags_0_io_debugSignals_20};
  assign regs_io_argOuts_23_bits = {{32'd0}, mags_0_io_debugSignals_21};
  assign regs_io_argOuts_24_bits = {{32'd0}, mags_0_io_debugSignals_22};
  assign regs_io_argOuts_25_bits = {{32'd0}, mags_0_io_debugSignals_23};
  assign regs_io_argOuts_26_bits = {{32'd0}, mags_0_io_debugSignals_24};
  assign regs_io_argOuts_27_bits = {{32'd0}, mags_0_io_debugSignals_25};
  assign regs_io_argOuts_28_bits = {{32'd0}, mags_0_io_debugSignals_26};
  assign regs_io_argOuts_29_bits = {{32'd0}, mags_0_io_debugSignals_27};
  assign regs_io_argOuts_30_bits = {{32'd0}, mags_0_io_debugSignals_28};
  assign regs_io_argOuts_31_bits = {{32'd0}, mags_0_io_debugSignals_29};
  assign regs_io_argOuts_32_bits = {{32'd0}, mags_0_io_debugSignals_30};
  assign regs_io_argOuts_33_bits = {{32'd0}, mags_0_io_debugSignals_31};
  assign regs_io_argOuts_34_bits = {{32'd0}, mags_0_io_debugSignals_32};
  assign regs_io_argOuts_35_bits = {{32'd0}, mags_0_io_debugSignals_33};
  assign regs_io_argOuts_36_bits = {{32'd0}, mags_0_io_debugSignals_34};
  assign regs_io_argOuts_37_bits = {{32'd0}, mags_0_io_debugSignals_35};
  assign regs_io_argOuts_38_bits = {{32'd0}, mags_0_io_debugSignals_36};
  assign regs_io_argOuts_39_bits = {{32'd0}, mags_0_io_debugSignals_37};
  assign regs_io_argOuts_40_bits = {{32'd0}, mags_0_io_debugSignals_38};
  assign regs_io_argOuts_41_bits = {{32'd0}, mags_0_io_debugSignals_39};
  assign regs_io_argOuts_42_bits = {{32'd0}, mags_0_io_debugSignals_40};
  assign regs_io_argOuts_43_bits = {{32'd0}, mags_0_io_debugSignals_41};
  assign regs_io_argOuts_44_bits = {{32'd0}, mags_0_io_debugSignals_42};
  assign regs_io_argOuts_45_bits = {{32'd0}, mags_0_io_debugSignals_43};
  assign regs_io_argOuts_46_bits = {{32'd0}, mags_0_io_debugSignals_44};
  assign regs_io_argOuts_47_bits = {{32'd0}, mags_0_io_debugSignals_45};
  assign regs_io_argOuts_48_bits = {{32'd0}, mags_0_io_debugSignals_46};
  assign regs_io_argOuts_49_bits = {{32'd0}, mags_0_io_debugSignals_47};
  assign regs_io_argOuts_50_bits = {{32'd0}, mags_0_io_debugSignals_48};
  assign regs_io_argOuts_51_bits = {{32'd0}, mags_0_io_debugSignals_49};
  assign regs_io_argOuts_52_bits = {{32'd0}, mags_0_io_debugSignals_50};
  assign regs_io_argOuts_53_bits = {{32'd0}, mags_0_io_debugSignals_51};
  assign regs_io_argOuts_54_bits = {{32'd0}, mags_0_io_debugSignals_52};
  assign regs_io_argOuts_55_bits = {{32'd0}, mags_0_io_debugSignals_53};
  assign regs_io_argOuts_56_bits = {{32'd0}, mags_0_io_debugSignals_54};
  assign regs_io_argOuts_57_bits = {{32'd0}, mags_0_io_debugSignals_55};
  assign regs_io_argOuts_58_bits = {{32'd0}, mags_0_io_debugSignals_56};
  assign regs_io_argOuts_59_bits = {{32'd0}, mags_0_io_debugSignals_57};
  assign regs_io_argOuts_60_bits = {{32'd0}, mags_0_io_debugSignals_58};
  assign regs_io_argOuts_61_bits = {{32'd0}, mags_0_io_debugSignals_59};
  assign regs_io_argOuts_62_bits = {{32'd0}, mags_0_io_debugSignals_60};
  assign regs_io_argOuts_63_bits = {{32'd0}, mags_0_io_debugSignals_61};
  assign regs_io_argOuts_64_bits = {{32'd0}, mags_0_io_debugSignals_62};
  assign regs_io_argOuts_65_bits = {{32'd0}, mags_0_io_debugSignals_63};
  assign regs_io_argOuts_66_bits = {{32'd0}, mags_0_io_debugSignals_64};
  assign regs_io_argOuts_67_bits = {{32'd0}, mags_0_io_debugSignals_65};
  assign regs_io_argOuts_68_bits = {{32'd0}, mags_0_io_debugSignals_66};
  assign regs_io_argOuts_69_bits = {{32'd0}, mags_0_io_debugSignals_67};
  assign regs_io_argOuts_70_bits = {{32'd0}, mags_0_io_debugSignals_68};
  assign regs_io_argOuts_71_bits = {{32'd0}, mags_0_io_debugSignals_69};
  assign regs_io_argOuts_72_bits = {{32'd0}, mags_0_io_debugSignals_70};
  assign regs_io_argOuts_73_bits = {{32'd0}, mags_0_io_debugSignals_71};
  assign regs_io_argOuts_74_bits = {{32'd0}, mags_0_io_debugSignals_72};
  assign regs_io_argOuts_75_bits = {{32'd0}, mags_0_io_debugSignals_73};
  assign regs_io_argOuts_76_bits = {{32'd0}, mags_0_io_debugSignals_74};
  assign regs_io_argOuts_77_bits = {{32'd0}, mags_0_io_debugSignals_75};
  assign regs_io_argOuts_78_bits = {{32'd0}, mags_0_io_debugSignals_76};
  assign regs_io_argOuts_79_bits = {{32'd0}, mags_0_io_debugSignals_77};
  assign regs_io_argOuts_80_bits = {{32'd0}, mags_0_io_debugSignals_78};
  assign regs_io_argOuts_81_bits = {{32'd0}, mags_0_io_debugSignals_79};
  assign regs_io_argOuts_82_bits = {{32'd0}, mags_0_io_debugSignals_80};
  assign regs_io_argOuts_83_bits = {{32'd0}, mags_0_io_debugSignals_81};
  assign regs_io_argOuts_84_bits = {{32'd0}, mags_0_io_debugSignals_82};
  assign regs_io_argOuts_85_bits = {{32'd0}, mags_0_io_debugSignals_83};
  assign regs_io_argOuts_86_bits = {{32'd0}, mags_0_io_debugSignals_84};
  assign regs_io_argOuts_87_bits = {{32'd0}, mags_0_io_debugSignals_85};
  assign regs_io_argOuts_88_bits = {{32'd0}, mags_0_io_debugSignals_86};
  assign regs_io_argOuts_89_bits = {{32'd0}, mags_0_io_debugSignals_87};
  assign regs_io_argOuts_90_bits = {{32'd0}, mags_0_io_debugSignals_88};
  assign regs_io_argOuts_91_bits = {{32'd0}, mags_0_io_debugSignals_89};
  assign regs_io_argOuts_92_bits = {{32'd0}, mags_0_io_debugSignals_90};
  assign regs_io_argOuts_93_bits = {{32'd0}, mags_0_io_debugSignals_91};
  assign regs_io_argOuts_94_bits = {{32'd0}, mags_0_io_debugSignals_92};
  assign regs_io_argOuts_95_bits = {{32'd0}, mags_0_io_debugSignals_93};
  assign regs_io_argOuts_96_bits = {{32'd0}, mags_0_io_debugSignals_94};
  assign regs_io_argOuts_97_bits = {{32'd0}, mags_0_io_debugSignals_95};
  assign regs_io_argOuts_98_bits = {{32'd0}, mags_0_io_debugSignals_96};
  assign regs_io_argOuts_99_bits = {{32'd0}, mags_0_io_debugSignals_97};
  assign regs_io_argOuts_100_bits = {{32'd0}, mags_0_io_debugSignals_98};
  assign regs_io_argOuts_101_bits = {{32'd0}, mags_0_io_debugSignals_99};
  assign regs_io_argOuts_102_bits = {{32'd0}, mags_0_io_debugSignals_100};
  assign regs_io_argOuts_103_bits = {{32'd0}, mags_0_io_debugSignals_101};
  assign regs_io_argOuts_104_bits = {{32'd0}, mags_0_io_debugSignals_102};
  assign regs_io_argOuts_105_bits = {{32'd0}, mags_0_io_debugSignals_103};
  assign regs_io_argOuts_106_bits = {{32'd0}, mags_0_io_debugSignals_104};
  assign regs_io_argOuts_107_bits = {{32'd0}, mags_0_io_debugSignals_105};
  assign regs_io_argOuts_108_bits = {{32'd0}, mags_0_io_debugSignals_106};
  assign regs_io_argOuts_109_bits = {{32'd0}, mags_0_io_debugSignals_107};
  assign regs_io_argOuts_110_bits = {{32'd0}, mags_0_io_debugSignals_108};
  assign regs_io_argOuts_111_bits = {{32'd0}, mags_0_io_debugSignals_109};
  assign regs_io_argOuts_112_bits = {{32'd0}, mags_0_io_debugSignals_110};
  assign regs_io_argOuts_113_bits = {{32'd0}, mags_0_io_debugSignals_111};
  assign regs_io_argOuts_114_bits = {{32'd0}, mags_0_io_debugSignals_112};
  assign regs_io_argOuts_115_bits = {{32'd0}, mags_0_io_debugSignals_113};
  assign regs_clock = clock;
  assign regs_reset = reset;
  assign timeoutCtr_io_enable = localEnable;
  assign timeoutCtr_clock = clock;
  assign timeoutCtr_reset = reset;
  assign depulser_io_in = _T_532;
  assign depulser_io_rst = _T_533[0];
  assign depulser_clock = clock;
  assign depulser_reset = reset;
  assign status_valid = depulser_io_out;
  assign status_bits = {{62'd0}, _T_546};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{$random}};
  _T_524 = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_524 <= _GEN_0;
  end
endmodule
module MAGToAXI4Bridge(
  output         io_in_cmd_ready,
  input          io_in_cmd_valid,
  input  [63:0]  io_in_cmd_bits_addr,
  input  [31:0]  io_in_cmd_bits_size,
  input          io_in_cmd_bits_isWr,
  input  [25:0]  io_in_cmd_bits_tag_uid,
  input  [5:0]   io_in_cmd_bits_tag_streamId,
  output         io_in_wdata_ready,
  input          io_in_wdata_valid,
  input  [31:0]  io_in_wdata_bits_wdata_0,
  input  [31:0]  io_in_wdata_bits_wdata_1,
  input  [31:0]  io_in_wdata_bits_wdata_2,
  input  [31:0]  io_in_wdata_bits_wdata_3,
  input  [31:0]  io_in_wdata_bits_wdata_4,
  input  [31:0]  io_in_wdata_bits_wdata_5,
  input  [31:0]  io_in_wdata_bits_wdata_6,
  input  [31:0]  io_in_wdata_bits_wdata_7,
  input  [31:0]  io_in_wdata_bits_wdata_8,
  input  [31:0]  io_in_wdata_bits_wdata_9,
  input  [31:0]  io_in_wdata_bits_wdata_10,
  input  [31:0]  io_in_wdata_bits_wdata_11,
  input  [31:0]  io_in_wdata_bits_wdata_12,
  input  [31:0]  io_in_wdata_bits_wdata_13,
  input  [31:0]  io_in_wdata_bits_wdata_14,
  input  [31:0]  io_in_wdata_bits_wdata_15,
  input          io_in_wdata_bits_wlast,
  input          io_in_rresp_ready,
  output         io_in_rresp_valid,
  output [31:0]  io_in_rresp_bits_rdata_0,
  output [31:0]  io_in_rresp_bits_rdata_1,
  output [31:0]  io_in_rresp_bits_rdata_2,
  output [31:0]  io_in_rresp_bits_rdata_3,
  output [31:0]  io_in_rresp_bits_rdata_4,
  output [31:0]  io_in_rresp_bits_rdata_5,
  output [31:0]  io_in_rresp_bits_rdata_6,
  output [31:0]  io_in_rresp_bits_rdata_7,
  output [31:0]  io_in_rresp_bits_rdata_8,
  output [31:0]  io_in_rresp_bits_rdata_9,
  output [31:0]  io_in_rresp_bits_rdata_10,
  output [31:0]  io_in_rresp_bits_rdata_11,
  output [31:0]  io_in_rresp_bits_rdata_12,
  output [31:0]  io_in_rresp_bits_rdata_13,
  output [31:0]  io_in_rresp_bits_rdata_14,
  output [31:0]  io_in_rresp_bits_rdata_15,
  output [5:0]   io_in_rresp_bits_tag_streamId,
  input          io_in_wresp_ready,
  output         io_in_wresp_valid,
  output [5:0]   io_in_wresp_bits_tag_streamId,
  output [5:0]   io_M_AXI_AWID,
  output [31:0]  io_M_AXI_AWADDR,
  output [7:0]   io_M_AXI_AWLEN,
  output         io_M_AXI_AWVALID,
  input          io_M_AXI_AWREADY,
  output [5:0]   io_M_AXI_ARID,
  output [31:0]  io_M_AXI_ARADDR,
  output [7:0]   io_M_AXI_ARLEN,
  output         io_M_AXI_ARVALID,
  input          io_M_AXI_ARREADY,
  output [511:0] io_M_AXI_WDATA,
  output         io_M_AXI_WLAST,
  output         io_M_AXI_WVALID,
  input          io_M_AXI_WREADY,
  input  [5:0]   io_M_AXI_RID,
  input  [511:0] io_M_AXI_RDATA,
  input          io_M_AXI_RVALID,
  output         io_M_AXI_RREADY,
  input  [5:0]   io_M_AXI_BID,
  input          io_M_AXI_BVALID,
  output         io_M_AXI_BREADY
);
  wire [31:0] id;
  wire [32:0] _T_125;
  wire [32:0] _T_126;
  wire [31:0] _T_127;
  wire  _T_134;
  wire  _T_135;
  wire  _T_136;
  wire  _T_147;
  wire [63:0] _T_148;
  wire [95:0] _T_149;
  wire [127:0] _T_150;
  wire [159:0] _T_151;
  wire [191:0] _T_152;
  wire [223:0] _T_153;
  wire [255:0] _T_154;
  wire [287:0] _T_155;
  wire [319:0] _T_156;
  wire [351:0] _T_157;
  wire [383:0] _T_158;
  wire [415:0] _T_159;
  wire [447:0] _T_160;
  wire [479:0] _T_161;
  wire [511:0] _T_162;
  wire [31:0] _T_168;
  wire [31:0] _T_169;
  wire [31:0] _T_170;
  wire [31:0] _T_171;
  wire [31:0] _T_172;
  wire [31:0] _T_173;
  wire [31:0] _T_174;
  wire [31:0] _T_175;
  wire [31:0] _T_176;
  wire [31:0] _T_177;
  wire [31:0] _T_178;
  wire [31:0] _T_179;
  wire [31:0] _T_180;
  wire [31:0] _T_181;
  wire [31:0] _T_182;
  wire [31:0] _T_183;
  wire [31:0] rdataAsVec_0;
  wire [31:0] rdataAsVec_1;
  wire [31:0] rdataAsVec_2;
  wire [31:0] rdataAsVec_3;
  wire [31:0] rdataAsVec_4;
  wire [31:0] rdataAsVec_5;
  wire [31:0] rdataAsVec_6;
  wire [31:0] rdataAsVec_7;
  wire [31:0] rdataAsVec_8;
  wire [31:0] rdataAsVec_9;
  wire [31:0] rdataAsVec_10;
  wire [31:0] rdataAsVec_11;
  wire [31:0] rdataAsVec_12;
  wire [31:0] rdataAsVec_13;
  wire [31:0] rdataAsVec_14;
  wire [31:0] rdataAsVec_15;
  wire [5:0] _T_206_streamId;
  wire [31:0] _T_208;
  wire [5:0] _T_209;
  wire [5:0] _T_213_streamId;
  wire [31:0] _T_215;
  wire [5:0] _T_216;
  assign id = {io_in_cmd_bits_tag_uid,io_in_cmd_bits_tag_streamId};
  assign _T_125 = io_in_cmd_bits_size - 32'h1;
  assign _T_126 = $unsigned(_T_125);
  assign _T_127 = _T_126[31:0];
  assign _T_134 = ~ io_in_cmd_bits_isWr;
  assign _T_135 = io_in_cmd_valid & _T_134;
  assign _T_136 = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY;
  assign _T_147 = io_in_cmd_valid & io_in_cmd_bits_isWr;
  assign _T_148 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14};
  assign _T_149 = {_T_148,io_in_wdata_bits_wdata_13};
  assign _T_150 = {_T_149,io_in_wdata_bits_wdata_12};
  assign _T_151 = {_T_150,io_in_wdata_bits_wdata_11};
  assign _T_152 = {_T_151,io_in_wdata_bits_wdata_10};
  assign _T_153 = {_T_152,io_in_wdata_bits_wdata_9};
  assign _T_154 = {_T_153,io_in_wdata_bits_wdata_8};
  assign _T_155 = {_T_154,io_in_wdata_bits_wdata_7};
  assign _T_156 = {_T_155,io_in_wdata_bits_wdata_6};
  assign _T_157 = {_T_156,io_in_wdata_bits_wdata_5};
  assign _T_158 = {_T_157,io_in_wdata_bits_wdata_4};
  assign _T_159 = {_T_158,io_in_wdata_bits_wdata_3};
  assign _T_160 = {_T_159,io_in_wdata_bits_wdata_2};
  assign _T_161 = {_T_160,io_in_wdata_bits_wdata_1};
  assign _T_162 = {_T_161,io_in_wdata_bits_wdata_0};
  assign _T_168 = io_M_AXI_RDATA[511:480];
  assign _T_169 = io_M_AXI_RDATA[479:448];
  assign _T_170 = io_M_AXI_RDATA[447:416];
  assign _T_171 = io_M_AXI_RDATA[415:384];
  assign _T_172 = io_M_AXI_RDATA[383:352];
  assign _T_173 = io_M_AXI_RDATA[351:320];
  assign _T_174 = io_M_AXI_RDATA[319:288];
  assign _T_175 = io_M_AXI_RDATA[287:256];
  assign _T_176 = io_M_AXI_RDATA[255:224];
  assign _T_177 = io_M_AXI_RDATA[223:192];
  assign _T_178 = io_M_AXI_RDATA[191:160];
  assign _T_179 = io_M_AXI_RDATA[159:128];
  assign _T_180 = io_M_AXI_RDATA[127:96];
  assign _T_181 = io_M_AXI_RDATA[95:64];
  assign _T_182 = io_M_AXI_RDATA[63:32];
  assign _T_183 = io_M_AXI_RDATA[31:0];
  assign _T_209 = _T_208[5:0];
  assign _T_216 = _T_215[5:0];
  assign io_in_cmd_ready = _T_136;
  assign io_in_wdata_ready = io_M_AXI_WREADY;
  assign io_in_rresp_valid = io_M_AXI_RVALID;
  assign io_in_rresp_bits_rdata_0 = rdataAsVec_0;
  assign io_in_rresp_bits_rdata_1 = rdataAsVec_1;
  assign io_in_rresp_bits_rdata_2 = rdataAsVec_2;
  assign io_in_rresp_bits_rdata_3 = rdataAsVec_3;
  assign io_in_rresp_bits_rdata_4 = rdataAsVec_4;
  assign io_in_rresp_bits_rdata_5 = rdataAsVec_5;
  assign io_in_rresp_bits_rdata_6 = rdataAsVec_6;
  assign io_in_rresp_bits_rdata_7 = rdataAsVec_7;
  assign io_in_rresp_bits_rdata_8 = rdataAsVec_8;
  assign io_in_rresp_bits_rdata_9 = rdataAsVec_9;
  assign io_in_rresp_bits_rdata_10 = rdataAsVec_10;
  assign io_in_rresp_bits_rdata_11 = rdataAsVec_11;
  assign io_in_rresp_bits_rdata_12 = rdataAsVec_12;
  assign io_in_rresp_bits_rdata_13 = rdataAsVec_13;
  assign io_in_rresp_bits_rdata_14 = rdataAsVec_14;
  assign io_in_rresp_bits_rdata_15 = rdataAsVec_15;
  assign io_in_rresp_bits_tag_streamId = _T_206_streamId;
  assign io_in_wresp_valid = io_M_AXI_BVALID;
  assign io_in_wresp_bits_tag_streamId = _T_213_streamId;
  assign io_M_AXI_AWID = id[5:0];
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0];
  assign io_M_AXI_AWLEN = _T_127[7:0];
  assign io_M_AXI_AWVALID = _T_147;
  assign io_M_AXI_ARID = id[5:0];
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0];
  assign io_M_AXI_ARLEN = _T_127[7:0];
  assign io_M_AXI_ARVALID = _T_135;
  assign io_M_AXI_WDATA = _T_162;
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast;
  assign io_M_AXI_WVALID = io_in_wdata_valid;
  assign io_M_AXI_RREADY = io_in_rresp_ready;
  assign io_M_AXI_BREADY = io_in_wresp_ready;
  assign rdataAsVec_0 = _T_183;
  assign rdataAsVec_1 = _T_182;
  assign rdataAsVec_2 = _T_181;
  assign rdataAsVec_3 = _T_180;
  assign rdataAsVec_4 = _T_179;
  assign rdataAsVec_5 = _T_178;
  assign rdataAsVec_6 = _T_177;
  assign rdataAsVec_7 = _T_176;
  assign rdataAsVec_8 = _T_175;
  assign rdataAsVec_9 = _T_174;
  assign rdataAsVec_10 = _T_173;
  assign rdataAsVec_11 = _T_172;
  assign rdataAsVec_12 = _T_171;
  assign rdataAsVec_13 = _T_170;
  assign rdataAsVec_14 = _T_169;
  assign rdataAsVec_15 = _T_168;
  assign _T_206_streamId = _T_209;
  assign _T_208 = {{26'd0}, io_M_AXI_RID};
  assign _T_213_streamId = _T_216;
  assign _T_215 = {{26'd0}, io_M_AXI_BID};
endmodule
module FringeArria10(
  input          clock,
  input          reset,
  output [31:0]  io_S_AVALON_readdata,
  input  [6:0]   io_S_AVALON_address,
  input          io_S_AVALON_write,
  input  [31:0]  io_S_AVALON_writedata,
  output [5:0]   io_M_AXI_0_AWID,
  output [31:0]  io_M_AXI_0_AWADDR,
  output [7:0]   io_M_AXI_0_AWLEN,
  output         io_M_AXI_0_AWVALID,
  input          io_M_AXI_0_AWREADY,
  output [5:0]   io_M_AXI_0_ARID,
  output [31:0]  io_M_AXI_0_ARADDR,
  output [7:0]   io_M_AXI_0_ARLEN,
  output         io_M_AXI_0_ARVALID,
  input          io_M_AXI_0_ARREADY,
  output [511:0] io_M_AXI_0_WDATA,
  output         io_M_AXI_0_WLAST,
  output         io_M_AXI_0_WVALID,
  input          io_M_AXI_0_WREADY,
  input  [5:0]   io_M_AXI_0_RID,
  input  [511:0] io_M_AXI_0_RDATA,
  input          io_M_AXI_0_RVALID,
  output         io_M_AXI_0_RREADY,
  input  [5:0]   io_M_AXI_0_BID,
  input          io_M_AXI_0_BVALID,
  output         io_M_AXI_0_BREADY,
  output         io_enable,
  input          io_done,
  output [31:0]  io_argIns_0,
  output [31:0]  io_argIns_1,
  input          io_argOuts_0_valid,
  input  [31:0]  io_argOuts_0_bits
);
  wire  fringeCommon_clock;
  wire  fringeCommon_reset;
  wire [31:0] fringeCommon_io_raddr;
  wire  fringeCommon_io_wen;
  wire [31:0] fringeCommon_io_waddr;
  wire [63:0] fringeCommon_io_wdata;
  wire [63:0] fringeCommon_io_rdata;
  wire  fringeCommon_io_enable;
  wire  fringeCommon_io_done;
  wire [63:0] fringeCommon_io_argIns_0;
  wire [63:0] fringeCommon_io_argIns_1;
  wire  fringeCommon_io_argOuts_0_valid;
  wire [63:0] fringeCommon_io_argOuts_0_bits;
  wire  fringeCommon_io_dram_0_cmd_ready;
  wire  fringeCommon_io_dram_0_cmd_valid;
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr;
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size;
  wire  fringeCommon_io_dram_0_cmd_bits_isWr;
  wire [25:0] fringeCommon_io_dram_0_cmd_bits_tag_uid;
  wire [5:0] fringeCommon_io_dram_0_cmd_bits_tag_streamId;
  wire  fringeCommon_io_dram_0_wdata_ready;
  wire  fringeCommon_io_dram_0_wdata_valid;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15;
  wire  fringeCommon_io_dram_0_wdata_bits_wlast;
  wire  fringeCommon_io_dram_0_rresp_ready;
  wire  fringeCommon_io_dram_0_rresp_valid;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_0;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_1;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_2;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_3;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_4;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_5;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_6;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_7;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_8;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_9;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_10;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_11;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_12;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_13;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_14;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_15;
  wire [5:0] fringeCommon_io_dram_0_rresp_bits_tag_streamId;
  wire  fringeCommon_io_dram_0_wresp_ready;
  wire  fringeCommon_io_dram_0_wresp_valid;
  wire [5:0] fringeCommon_io_dram_0_wresp_bits_tag_streamId;
  wire  MAGToAXI4Bridge_io_in_cmd_ready;
  wire  MAGToAXI4Bridge_io_in_cmd_valid;
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr;
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size;
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr;
  wire [25:0] MAGToAXI4Bridge_io_in_cmd_bits_tag_uid;
  wire [5:0] MAGToAXI4Bridge_io_in_cmd_bits_tag_streamId;
  wire  MAGToAXI4Bridge_io_in_wdata_ready;
  wire  MAGToAXI4Bridge_io_in_wdata_valid;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast;
  wire  MAGToAXI4Bridge_io_in_rresp_ready;
  wire  MAGToAXI4Bridge_io_in_rresp_valid;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_0;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_1;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_2;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_3;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_4;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_5;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_6;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_7;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_8;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_9;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_10;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_11;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_12;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_13;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_14;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_15;
  wire [5:0] MAGToAXI4Bridge_io_in_rresp_bits_tag_streamId;
  wire  MAGToAXI4Bridge_io_in_wresp_ready;
  wire  MAGToAXI4Bridge_io_in_wresp_valid;
  wire [5:0] MAGToAXI4Bridge_io_in_wresp_bits_tag_streamId;
  wire [5:0] MAGToAXI4Bridge_io_M_AXI_AWID;
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR;
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN;
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID;
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY;
  wire [5:0] MAGToAXI4Bridge_io_M_AXI_ARID;
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR;
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN;
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID;
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY;
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA;
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST;
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID;
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY;
  wire [5:0] MAGToAXI4Bridge_io_M_AXI_RID;
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_RDATA;
  wire  MAGToAXI4Bridge_io_M_AXI_RVALID;
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY;
  wire [5:0] MAGToAXI4Bridge_io_M_AXI_BID;
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID;
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY;
  Fringe fringeCommon (
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag_uid(fringeCommon_io_dram_0_cmd_bits_tag_uid),
    .io_dram_0_cmd_bits_tag_streamId(fringeCommon_io_dram_0_cmd_bits_tag_streamId),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_rresp_valid(fringeCommon_io_dram_0_rresp_valid),
    .io_dram_0_rresp_bits_rdata_0(fringeCommon_io_dram_0_rresp_bits_rdata_0),
    .io_dram_0_rresp_bits_rdata_1(fringeCommon_io_dram_0_rresp_bits_rdata_1),
    .io_dram_0_rresp_bits_rdata_2(fringeCommon_io_dram_0_rresp_bits_rdata_2),
    .io_dram_0_rresp_bits_rdata_3(fringeCommon_io_dram_0_rresp_bits_rdata_3),
    .io_dram_0_rresp_bits_rdata_4(fringeCommon_io_dram_0_rresp_bits_rdata_4),
    .io_dram_0_rresp_bits_rdata_5(fringeCommon_io_dram_0_rresp_bits_rdata_5),
    .io_dram_0_rresp_bits_rdata_6(fringeCommon_io_dram_0_rresp_bits_rdata_6),
    .io_dram_0_rresp_bits_rdata_7(fringeCommon_io_dram_0_rresp_bits_rdata_7),
    .io_dram_0_rresp_bits_rdata_8(fringeCommon_io_dram_0_rresp_bits_rdata_8),
    .io_dram_0_rresp_bits_rdata_9(fringeCommon_io_dram_0_rresp_bits_rdata_9),
    .io_dram_0_rresp_bits_rdata_10(fringeCommon_io_dram_0_rresp_bits_rdata_10),
    .io_dram_0_rresp_bits_rdata_11(fringeCommon_io_dram_0_rresp_bits_rdata_11),
    .io_dram_0_rresp_bits_rdata_12(fringeCommon_io_dram_0_rresp_bits_rdata_12),
    .io_dram_0_rresp_bits_rdata_13(fringeCommon_io_dram_0_rresp_bits_rdata_13),
    .io_dram_0_rresp_bits_rdata_14(fringeCommon_io_dram_0_rresp_bits_rdata_14),
    .io_dram_0_rresp_bits_rdata_15(fringeCommon_io_dram_0_rresp_bits_rdata_15),
    .io_dram_0_rresp_bits_tag_streamId(fringeCommon_io_dram_0_rresp_bits_tag_streamId),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag_streamId(fringeCommon_io_dram_0_wresp_bits_tag_streamId)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge (
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag_uid(MAGToAXI4Bridge_io_in_cmd_bits_tag_uid),
    .io_in_cmd_bits_tag_streamId(MAGToAXI4Bridge_io_in_cmd_bits_tag_streamId),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_rresp_valid(MAGToAXI4Bridge_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(MAGToAXI4Bridge_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(MAGToAXI4Bridge_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(MAGToAXI4Bridge_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(MAGToAXI4Bridge_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(MAGToAXI4Bridge_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(MAGToAXI4Bridge_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(MAGToAXI4Bridge_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(MAGToAXI4Bridge_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_rdata_8(MAGToAXI4Bridge_io_in_rresp_bits_rdata_8),
    .io_in_rresp_bits_rdata_9(MAGToAXI4Bridge_io_in_rresp_bits_rdata_9),
    .io_in_rresp_bits_rdata_10(MAGToAXI4Bridge_io_in_rresp_bits_rdata_10),
    .io_in_rresp_bits_rdata_11(MAGToAXI4Bridge_io_in_rresp_bits_rdata_11),
    .io_in_rresp_bits_rdata_12(MAGToAXI4Bridge_io_in_rresp_bits_rdata_12),
    .io_in_rresp_bits_rdata_13(MAGToAXI4Bridge_io_in_rresp_bits_rdata_13),
    .io_in_rresp_bits_rdata_14(MAGToAXI4Bridge_io_in_rresp_bits_rdata_14),
    .io_in_rresp_bits_rdata_15(MAGToAXI4Bridge_io_in_rresp_bits_rdata_15),
    .io_in_rresp_bits_tag_streamId(MAGToAXI4Bridge_io_in_rresp_bits_tag_streamId),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag_streamId(MAGToAXI4Bridge_io_in_wresp_bits_tag_streamId),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RID(MAGToAXI4Bridge_io_M_AXI_RID),
    .io_M_AXI_RDATA(MAGToAXI4Bridge_io_M_AXI_RDATA),
    .io_M_AXI_RVALID(MAGToAXI4Bridge_io_M_AXI_RVALID),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  assign io_S_AVALON_readdata = fringeCommon_io_rdata[31:0];
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID;
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR;
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN;
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID;
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID;
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR;
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN;
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID;
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA;
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST;
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID;
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY;
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY;
  assign io_enable = fringeCommon_io_enable;
  assign io_argIns_0 = fringeCommon_io_argIns_0[31:0];
  assign io_argIns_1 = fringeCommon_io_argIns_1[31:0];
  assign fringeCommon_io_raddr = {{25'd0}, io_S_AVALON_address};
  assign fringeCommon_io_wen = io_S_AVALON_write;
  assign fringeCommon_io_waddr = {{25'd0}, io_S_AVALON_address};
  assign fringeCommon_io_wdata = {{32'd0}, io_S_AVALON_writedata};
  assign fringeCommon_io_done = io_done;
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid;
  assign fringeCommon_io_argOuts_0_bits = {{32'd0}, io_argOuts_0_bits};
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready;
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready;
  assign fringeCommon_io_dram_0_rresp_valid = MAGToAXI4Bridge_io_in_rresp_valid;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_0 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_0;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_1 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_1;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_2 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_2;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_3 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_3;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_4 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_4;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_5 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_5;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_6 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_6;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_7 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_7;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_8 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_8;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_9 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_9;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_10 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_10;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_11 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_11;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_12 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_12;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_13 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_13;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_14 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_14;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_15 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_15;
  assign fringeCommon_io_dram_0_rresp_bits_tag_streamId = MAGToAXI4Bridge_io_in_rresp_bits_tag_streamId;
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid;
  assign fringeCommon_io_dram_0_wresp_bits_tag_streamId = MAGToAXI4Bridge_io_in_wresp_bits_tag_streamId;
  assign fringeCommon_clock = clock;
  assign fringeCommon_reset = reset;
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid;
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr;
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size;
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr;
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag_uid = fringeCommon_io_dram_0_cmd_bits_tag_uid;
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag_streamId = fringeCommon_io_dram_0_cmd_bits_tag_streamId;
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast;
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready;
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready;
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY;
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY;
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY;
  assign MAGToAXI4Bridge_io_M_AXI_RID = io_M_AXI_0_RID;
  assign MAGToAXI4Bridge_io_M_AXI_RDATA = io_M_AXI_0_RDATA;
  assign MAGToAXI4Bridge_io_M_AXI_RVALID = io_M_AXI_0_RVALID;
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID;
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID;
endmodule
module Top(
  input          clock,
  input          reset,
  input          io_raddr,
  input          io_wen,
  input          io_waddr,
  input          io_wdata,
  output         io_rdata,
  output         io_is_enabled,
  output [31:0]  io_S_AVALON_readdata,
  input  [6:0]   io_S_AVALON_address,
  input          io_S_AVALON_chipselect,
  input          io_S_AVALON_write,
  input          io_S_AVALON_read,
  input  [31:0]  io_S_AVALON_writedata,
  output [5:0]   io_M_AXI_0_AWID,
  output [31:0]  io_M_AXI_0_AWUSER,
  output [31:0]  io_M_AXI_0_AWADDR,
  output [7:0]   io_M_AXI_0_AWLEN,
  output [2:0]   io_M_AXI_0_AWSIZE,
  output [1:0]   io_M_AXI_0_AWBURST,
  output         io_M_AXI_0_AWLOCK,
  output [3:0]   io_M_AXI_0_AWCACHE,
  output [2:0]   io_M_AXI_0_AWPROT,
  output [3:0]   io_M_AXI_0_AWQOS,
  output         io_M_AXI_0_AWVALID,
  input          io_M_AXI_0_AWREADY,
  output [5:0]   io_M_AXI_0_ARID,
  output [31:0]  io_M_AXI_0_ARUSER,
  output [31:0]  io_M_AXI_0_ARADDR,
  output [7:0]   io_M_AXI_0_ARLEN,
  output [2:0]   io_M_AXI_0_ARSIZE,
  output [1:0]   io_M_AXI_0_ARBURST,
  output         io_M_AXI_0_ARLOCK,
  output [3:0]   io_M_AXI_0_ARCACHE,
  output [2:0]   io_M_AXI_0_ARPROT,
  output [3:0]   io_M_AXI_0_ARQOS,
  output         io_M_AXI_0_ARVALID,
  input          io_M_AXI_0_ARREADY,
  output [511:0] io_M_AXI_0_WDATA,
  output [63:0]  io_M_AXI_0_WSTRB,
  output         io_M_AXI_0_WLAST,
  output         io_M_AXI_0_WVALID,
  input          io_M_AXI_0_WREADY,
  input  [5:0]   io_M_AXI_0_RID,
  input  [31:0]  io_M_AXI_0_RUSER,
  input  [511:0] io_M_AXI_0_RDATA,
  input  [1:0]   io_M_AXI_0_RRESP,
  input          io_M_AXI_0_RLAST,
  input          io_M_AXI_0_RVALID,
  output         io_M_AXI_0_RREADY,
  input  [5:0]   io_M_AXI_0_BID,
  input  [31:0]  io_M_AXI_0_BUSER,
  input  [1:0]   io_M_AXI_0_BRESP,
  input          io_M_AXI_0_BVALID,
  output         io_M_AXI_0_BREADY
);
  wire  accel_clock;
  wire  accel_reset;
  wire  accel_io_enable;
  wire  accel_io_done;
  wire [63:0] accel_io_argIns_0;
  wire [63:0] accel_io_argIns_1;
  wire  accel_io_argOuts_0_valid;
  wire [63:0] accel_io_argOuts_0_bits;
  wire  FringeArria10_clock;
  wire  FringeArria10_reset;
  wire [31:0] FringeArria10_io_S_AVALON_readdata;
  wire [6:0] FringeArria10_io_S_AVALON_address;
  wire  FringeArria10_io_S_AVALON_write;
  wire [31:0] FringeArria10_io_S_AVALON_writedata;
  wire [5:0] FringeArria10_io_M_AXI_0_AWID;
  wire [31:0] FringeArria10_io_M_AXI_0_AWADDR;
  wire [7:0] FringeArria10_io_M_AXI_0_AWLEN;
  wire  FringeArria10_io_M_AXI_0_AWVALID;
  wire  FringeArria10_io_M_AXI_0_AWREADY;
  wire [5:0] FringeArria10_io_M_AXI_0_ARID;
  wire [31:0] FringeArria10_io_M_AXI_0_ARADDR;
  wire [7:0] FringeArria10_io_M_AXI_0_ARLEN;
  wire  FringeArria10_io_M_AXI_0_ARVALID;
  wire  FringeArria10_io_M_AXI_0_ARREADY;
  wire [511:0] FringeArria10_io_M_AXI_0_WDATA;
  wire  FringeArria10_io_M_AXI_0_WLAST;
  wire  FringeArria10_io_M_AXI_0_WVALID;
  wire  FringeArria10_io_M_AXI_0_WREADY;
  wire [5:0] FringeArria10_io_M_AXI_0_RID;
  wire [511:0] FringeArria10_io_M_AXI_0_RDATA;
  wire  FringeArria10_io_M_AXI_0_RVALID;
  wire  FringeArria10_io_M_AXI_0_RREADY;
  wire [5:0] FringeArria10_io_M_AXI_0_BID;
  wire  FringeArria10_io_M_AXI_0_BVALID;
  wire  FringeArria10_io_M_AXI_0_BREADY;
  wire  FringeArria10_io_enable;
  wire  FringeArria10_io_done;
  wire [31:0] FringeArria10_io_argIns_0;
  wire [31:0] FringeArria10_io_argIns_1;
  wire  FringeArria10_io_argOuts_0_valid;
  wire [31:0] FringeArria10_io_argOuts_0_bits;
  AccelTop accel (
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_valid(accel_io_argOuts_0_valid),
    .io_argOuts_0_bits(accel_io_argOuts_0_bits)
  );
  FringeArria10 FringeArria10 (
    .clock(FringeArria10_clock),
    .reset(FringeArria10_reset),
    .io_S_AVALON_readdata(FringeArria10_io_S_AVALON_readdata),
    .io_S_AVALON_address(FringeArria10_io_S_AVALON_address),
    .io_S_AVALON_write(FringeArria10_io_S_AVALON_write),
    .io_S_AVALON_writedata(FringeArria10_io_S_AVALON_writedata),
    .io_M_AXI_0_AWID(FringeArria10_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeArria10_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeArria10_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeArria10_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeArria10_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeArria10_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeArria10_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeArria10_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeArria10_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeArria10_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeArria10_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WLAST(FringeArria10_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeArria10_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeArria10_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RID(FringeArria10_io_M_AXI_0_RID),
    .io_M_AXI_0_RDATA(FringeArria10_io_M_AXI_0_RDATA),
    .io_M_AXI_0_RVALID(FringeArria10_io_M_AXI_0_RVALID),
    .io_M_AXI_0_RREADY(FringeArria10_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeArria10_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeArria10_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeArria10_io_M_AXI_0_BREADY),
    .io_enable(FringeArria10_io_enable),
    .io_done(FringeArria10_io_done),
    .io_argIns_0(FringeArria10_io_argIns_0),
    .io_argIns_1(FringeArria10_io_argIns_1),
    .io_argOuts_0_valid(FringeArria10_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeArria10_io_argOuts_0_bits)
  );
  assign io_rdata = 1'h0;
  assign io_is_enabled = 1'h0;
  assign io_S_AVALON_readdata = FringeArria10_io_S_AVALON_readdata;
  assign io_M_AXI_0_AWID = FringeArria10_io_M_AXI_0_AWID;
  assign io_M_AXI_0_AWUSER = 32'h0;
  assign io_M_AXI_0_AWADDR = FringeArria10_io_M_AXI_0_AWADDR;
  assign io_M_AXI_0_AWLEN = FringeArria10_io_M_AXI_0_AWLEN;
  assign io_M_AXI_0_AWSIZE = 3'h6;
  assign io_M_AXI_0_AWBURST = 2'h1;
  assign io_M_AXI_0_AWLOCK = 1'h0;
  assign io_M_AXI_0_AWCACHE = 4'h3;
  assign io_M_AXI_0_AWPROT = 3'h0;
  assign io_M_AXI_0_AWQOS = 4'h0;
  assign io_M_AXI_0_AWVALID = FringeArria10_io_M_AXI_0_AWVALID;
  assign io_M_AXI_0_ARID = FringeArria10_io_M_AXI_0_ARID;
  assign io_M_AXI_0_ARUSER = 32'h0;
  assign io_M_AXI_0_ARADDR = FringeArria10_io_M_AXI_0_ARADDR;
  assign io_M_AXI_0_ARLEN = FringeArria10_io_M_AXI_0_ARLEN;
  assign io_M_AXI_0_ARSIZE = 3'h6;
  assign io_M_AXI_0_ARBURST = 2'h1;
  assign io_M_AXI_0_ARLOCK = 1'h0;
  assign io_M_AXI_0_ARCACHE = 4'h3;
  assign io_M_AXI_0_ARPROT = 3'h0;
  assign io_M_AXI_0_ARQOS = 4'h0;
  assign io_M_AXI_0_ARVALID = FringeArria10_io_M_AXI_0_ARVALID;
  assign io_M_AXI_0_WDATA = FringeArria10_io_M_AXI_0_WDATA;
  assign io_M_AXI_0_WSTRB = 64'hffffffffffffffff;
  assign io_M_AXI_0_WLAST = FringeArria10_io_M_AXI_0_WLAST;
  assign io_M_AXI_0_WVALID = FringeArria10_io_M_AXI_0_WVALID;
  assign io_M_AXI_0_RREADY = FringeArria10_io_M_AXI_0_RREADY;
  assign io_M_AXI_0_BREADY = FringeArria10_io_M_AXI_0_BREADY;
  assign accel_io_enable = FringeArria10_io_enable;
  assign accel_io_argIns_0 = {{32'd0}, FringeArria10_io_argIns_0};
  assign accel_io_argIns_1 = {{32'd0}, FringeArria10_io_argIns_1};
  assign accel_clock = clock;
  assign accel_reset = reset;
  assign FringeArria10_io_S_AVALON_address = io_S_AVALON_address;
  assign FringeArria10_io_S_AVALON_write = io_S_AVALON_write;
  assign FringeArria10_io_S_AVALON_writedata = io_S_AVALON_writedata;
  assign FringeArria10_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY;
  assign FringeArria10_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY;
  assign FringeArria10_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY;
  assign FringeArria10_io_M_AXI_0_RID = io_M_AXI_0_RID;
  assign FringeArria10_io_M_AXI_0_RDATA = io_M_AXI_0_RDATA;
  assign FringeArria10_io_M_AXI_0_RVALID = io_M_AXI_0_RVALID;
  assign FringeArria10_io_M_AXI_0_BID = io_M_AXI_0_BID;
  assign FringeArria10_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID;
  assign FringeArria10_io_done = accel_io_done;
  assign FringeArria10_io_argOuts_0_valid = accel_io_argOuts_0_valid;
  assign FringeArria10_io_argOuts_0_bits = accel_io_argOuts_0_bits[31:0];
  assign FringeArria10_clock = clock;
  assign FringeArria10_reset = reset;
endmodule
